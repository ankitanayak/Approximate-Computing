library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
 
entity adder_approxadder is
   port
   (
	approx_flag : in std_logic;
	bit_op1 : in std_logic;
      	bit_op2 : in std_logic;
	bit_cin : in std_logic;
	bit_sum : out std_logic;
	bit_cout : out std_logic
   );
end entity adder_approxadder;

architecture behav_adder_approxadder of adder_approxadder is

begin
   	process (bit_op1, bit_op2, bit_cin, approx_flag) is
   	begin
		if bit_op1 = '0' and bit_op2 = '0' and bit_cin = '0' then
			bit_sum <= '0';
			bit_cout <= '0';
		elsif bit_op1 = '0' and bit_op2 = '0' and bit_cin = '1' and approx_flag = '0' then
			bit_sum <= '1';
			bit_cout <= '0';
		elsif bit_op1 = '0' and bit_op2 = '0' and bit_cin = '1' and approx_flag = '1' then
			bit_sum <= '0';
			bit_cout <= '0';
		elsif bit_op1 = '0' and bit_op2 = '1' and bit_cin = '0' then
			bit_sum <= '1';
			bit_cout <= '0';
		elsif bit_op1 = '0' and bit_op2 = '1' and bit_cin = '1' and approx_flag = '0' then
			bit_sum <= '0';
			bit_cout <= '1';
		elsif bit_op1 = '0' and bit_op2 = '1' and bit_cin = '1' and approx_flag = '1' then
			bit_sum <= '1';
			bit_cout <= '0';
		elsif bit_op1 = '1' and bit_op2 = '0' and bit_cin = '0' and approx_flag = '0' then
			bit_sum <= '1';
			bit_cout <= '0';
		elsif bit_op1 = '1' and bit_op2 = '0' and bit_cin = '0' and approx_flag = '1' then
			bit_sum <= '0';
			bit_cout <= '1';
		elsif bit_op1 = '1' and bit_op2 = '0' and bit_cin = '1' then
			bit_sum <= '0';
			bit_cout <= '1';
		elsif bit_op1 = '1' and bit_op2 = '1' and bit_cin = '0' and approx_flag = '0' then
			bit_sum <= '0';
			bit_cout <= '1';
		elsif bit_op1 = '1' and bit_op2 = '1' and bit_cin = '0' and approx_flag = '1' then
			bit_sum <= '1';
			bit_cout <= '1';
		elsif bit_op1 = '1' and bit_op2 = '1' and bit_cin = '1' then
			bit_sum <= '1';
			bit_cout <= '1';
		end if;
	end process;
end architecture behav_adder_approxadder;
