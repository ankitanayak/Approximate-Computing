library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use IEEE.STD_LOGIC_TEXTIO.ALL;
use STD.TEXTIO.ALL;

entity blur is
   port
   (
	blur_xnor_value : in std_logic_vector (12 downto 0);
	blur_out_flag : out std_logic
   );
end entity blur;

architecture blur_arch of blur is

component blur_mult
port
   (
	blur_mult_regxnor_value : in std_logic_vector (12 downto 0);
	blur_mult_regop1 : in std_logic_vector (11 downto 0);
      	blur_mult_regop2 : in std_logic_vector (11 downto 0);
	blur_mult_regres : out std_logic_vector (23 downto 0)
   );
end component;

constant key_width: integer:=13;
constant matrix_size: integer:=128;
constant operand_width: integer:=12;
constant result_width: integer:=operand_width*2;

type blur_matrix_row_type is array (0 to matrix_size-1) of integer;
type blur_matrix_type is array (0 to matrix_size-1) of blur_matrix_row_type;

type blur_sum_matrix_row_type is array (0 to matrix_size-1) of std_logic_vector(operand_width-1 downto 0);
type blur_sum_matrix_type is array (0 to matrix_size-1) of blur_sum_matrix_row_type;

type blur_res_matrix_row_type is array (0 to matrix_size-1) of std_logic_vector(result_width-1 downto 0);
type blur_res_matrix_type is array (0 to matrix_size-1) of blur_res_matrix_row_type;

type blur_matrix_int_type is array (0 to (matrix_size*matrix_size)-1) of integer;

signal blur_matrix : blur_matrix_type;
signal blur_sum_matrix : blur_sum_matrix_type;
signal blur_res_matrix : blur_res_matrix_type;
signal blur_matrix_int : blur_matrix_int_type;

begin

	blur_matrix_int <=(137,135,136,133,135,130,129,129,131,137,144,151,149,138,118,86,62,65,72,74,76,77,76,77,77,75,80,85,87,92,93,96,100,98,103,98,97,101,99,103,100,103,101,101,103,101,102,102,104,105,104,104,105,101,101,100,103,103,98,99,104,104,101,102,107,98,100,101,99,101,99,99,98,97,97,98,91,90,86,75,79,102,117,129,137,136,123,127,128,129,131,128,126,126,128,129,131,132,135,129,141,192,208,213,209,137,72,78,89,93,93,90,94,92,89,90,92,95,95,90,96,96,95,93,84,89,139,136,
134,132,134,129,130,128,127,129,129,136,145,149,149,138,113,83,60,61,66,74,73,73,72,74,74,74,79,85,88,93,92,93,98,98,100,98,98,99,97,100,100,101,101,102,101,99,101,100,102,101,102,101,103,102,99,98,102,103,97,100,101,102,98,101,103,99,97,97,97,98,97,98,97,96,95,95,92,88,84,75,77,98,116,128,138,133,126,126,126,128,129,128,127,126,129,128,130,130,133,129,133,181,207,213,212,161,77,76,86,89,92,91,94,92,91,92,95,94,94,92,94,95,96,94,88,96,101,73,
132,129,132,129,129,130,126,127,129,140,145,148,148,133,109,82,57,55,64,69,70,70,73,71,70,74,79,83,87,92,91,94,94,96,97,98,100,98,98,99,99,102,100,99,100,99,100,99,99,99,100,97,99,100,98,96,100,99,96,98,100,99,97,97,99,99,97,96,96,96,94,95,96,96,96,95,92,88,83,77,73,84,106,120,131,135,130,127,131,131,131,131,130,128,129,127,129,128,128,129,125,147,196,209,214,202,121,70,81,86,90,92,91,92,90,92,94,92,92,92,93,94,93,102,101,72,29,16,
131,130,131,130,129,128,126,129,137,144,147,146,144,131,106,80,59,57,64,68,72,76,73,69,69,72,79,82,86,91,92,94,94,95,96,99,99,96,98,97,99,99,99,101,100,98,100,98,98,99,98,98,100,99,98,97,97,98,97,99,102,101,100,99,98,100,99,97,97,96,96,97,95,96,97,96,93,90,84,83,76,75,97,116,125,135,136,133,133,136,138,134,131,130,130,128,128,127,125,129,126,124,171,204,214,215,177,89,74,82,86,89,91,91,89,91,92,91,93,93,94,96,100,102,69,30,20,23,
130,129,130,131,131,128,127,133,142,145,143,143,139,126,108,83,58,58,64,68,73,73,70,71,70,69,78,82,86,89,93,93,95,96,96,98,98,98,99,97,99,98,98,102,100,99,99,99,96,101,100,99,100,100,100,97,99,101,96,98,102,105,101,99,100,99,98,95,98,97,95,93,96,98,96,97,94,91,85,83,78,72,86,110,122,130,138,138,135,138,140,136,134,133,131,127,128,126,126,126,125,121,138,192,211,215,210,142,72,78,85,86,91,92,92,94,93,96,96,96,98,103,103,63,22,20,22,22,
130,129,131,133,133,129,128,135,144,142,142,139,136,129,110,88,61,58,64,69,73,70,71,70,71,71,78,81,86,88,89,91,95,96,97,97,98,99,98,97,98,99,97,98,97,96,96,99,98,97,96,98,96,95,98,98,99,98,95,97,100,104,103,99,98,98,98,95,97,95,93,93,94,96,92,95,93,93,90,80,79,74,81,103,122,130,139,138,137,136,137,138,136,131,130,129,127,126,126,126,126,123,118,161,204,212,217,191,102,74,82,87,87,91,93,92,92,98,98,100,105,106,63,25,23,26,22,25,
129,129,131,132,132,129,132,140,145,142,139,135,135,130,109,79,57,55,62,70,71,71,73,70,69,72,76,80,87,89,89,93,96,94,95,96,96,95,96,98,97,96,95,98,96,94,96,99,103,97,92,92,90,91,93,94,93,92,94,94,96,97,100,98,99,99,96,94,94,94,93,94,95,93,93,95,92,92,92,79,77,74,84,99,118,130,136,138,137,135,135,135,136,133,131,130,128,127,125,126,126,123,118,129,187,210,215,216,159,76,79,88,92,92,93,90,89,93,97,102,106,60,29,20,19,20,23,26,
131,132,131,133,134,134,140,146,146,140,134,133,137,132,109,80,56,55,63,68,73,73,73,70,70,71,74,81,86,90,90,94,95,94,95,95,93,97,98,96,97,98,96,97,96,95,94,98,102,99,93,90,88,88,91,95,92,93,90,93,95,97,97,98,99,99,94,95,94,96,94,93,93,91,94,95,94,88,87,83,77,74,83,100,113,128,133,135,136,133,134,134,134,132,129,130,128,129,131,128,126,125,121,114,152,203,213,219,206,119,73,83,88,90,93,91,92,93,101,103,58,16,17,20,21,21,22,30,
132,133,135,135,136,140,146,146,144,139,133,133,136,131,109,80,57,59,64,66,72,73,72,68,68,70,76,80,83,88,90,91,93,94,94,95,93,92,93,96,95,95,97,96,96,97,95,96,98,95,93,89,89,87,88,92,94,91,90,91,93,96,97,97,101,98,95,95,96,94,94,92,93,93,92,95,94,88,85,82,78,73,83,96,109,121,129,133,135,133,132,135,132,132,132,131,130,128,130,130,128,126,123,116,119,179,210,218,221,183,89,73,83,86,92,93,95,100,103,61,18,15,27,25,25,23,25,26,
134,134,138,136,141,145,144,142,141,135,132,135,136,129,107,79,53,54,64,68,69,70,69,70,69,71,75,80,85,86,87,90,91,94,93,94,91,90,91,94,94,93,93,95,97,97,94,93,95,92,90,90,91,88,90,90,90,86,87,89,91,95,95,100,98,98,94,94,95,94,93,91,92,91,93,93,91,87,84,85,81,73,80,95,106,119,127,128,131,131,132,132,131,130,131,128,131,131,129,128,127,124,122,119,110,141,201,217,220,215,141,67,77,82,88,92,101,101,59,18,14,21,30,32,27,23,23,21,
135,136,136,138,145,142,136,135,135,135,132,135,136,128,107,77,51,53,63,70,69,68,70,69,68,70,74,80,86,87,88,91,90,89,92,92,90,90,94,93,93,92,93,94,94,94,94,93,94,93,92,93,87,88,85,85,85,85,82,80,83,90,94,97,98,93,93,92,93,97,91,93,93,92,93,92,91,88,83,83,81,76,80,92,107,115,121,127,128,131,131,128,129,129,128,126,128,130,127,125,123,120,118,116,112,114,176,214,219,222,195,96,69,79,82,93,100,62,19,16,20,26,32,29,26,22,19,19,
137,136,135,143,145,133,125,125,127,138,135,134,137,129,109,80,53,53,62,68,70,72,71,70,69,71,76,80,85,87,89,91,91,92,92,91,91,95,94,94,93,91,96,95,97,93,92,91,95,91,91,97,103,101,109,134,141,137,136,125,107,91,83,85,89,90,92,94,94,99,95,92,93,92,92,94,92,88,84,81,80,73,78,89,104,114,118,119,124,129,129,129,126,127,126,128,127,126,124,121,120,118,115,114,115,110,136,198,215,221,217,152,74,78,86,95,60,20,18,19,22,30,35,30,25,20,20,20,
135,134,136,148,140,123,116,113,123,139,137,135,138,129,109,81,54,54,59,65,70,71,69,70,69,71,77,79,84,87,88,91,93,91,92,92,94,93,95,94,94,92,93,96,97,92,91,90,103,116,119,126,126,142,150,159,168,168,172,175,169,165,139,110,86,82,87,91,98,97,97,93,92,91,90,92,88,85,85,79,78,73,75,91,104,116,114,118,121,124,128,128,125,125,127,126,126,123,121,118,116,114,112,112,112,111,113,163,209,216,222,204,114,78,92,61,15,15,18,20,27,29,32,30,20,16,18,20,
133,136,143,146,132,114,101,104,124,139,138,137,139,130,109,78,50,52,58,64,68,69,70,69,70,71,78,81,85,87,88,90,92,91,89,95,95,93,93,94,93,90,90,92,94,93,95,115,121,130,122,123,132,148,149,155,165,169,162,158,169,175,182,182,165,118,80,81,90,94,93,93,91,92,90,90,86,84,82,79,80,74,76,92,106,115,115,114,118,120,126,125,125,123,124,121,121,120,116,114,114,110,110,111,114,111,109,123,189,215,222,224,182,99,63,18,14,21,22,26,30,26,23,23,25,22,19,18,
134,139,149,138,121,98,83,105,129,142,141,139,139,132,111,76,47,47,59,62,65,66,67,66,70,71,76,81,83,85,88,88,89,88,89,92,91,92,94,91,89,95,106,114,109,94,106,118,118,117,122,128,125,134,141,149,154,160,162,164,165,173,176,182,191,189,154,93,78,89,92,91,87,90,89,87,85,82,78,79,75,74,78,89,107,115,117,115,116,118,121,124,124,120,118,118,116,117,115,112,112,110,109,109,109,111,110,106,146,208,218,225,226,127,15,13,19,21,28,27,26,27,22,24,26,21,21,21,
138,148,145,129,107,72,72,107,131,142,142,140,139,132,112,77,48,48,56,61,66,64,66,67,68,71,74,78,83,83,88,86,87,88,88,90,90,91,89,94,99,117,117,108,95,91,98,110,106,106,114,119,130,131,142,145,151,154,162,168,174,174,176,181,182,186,195,179,122,81,77,86,88,87,84,86,84,82,78,76,73,68,74,88,106,116,117,115,114,118,117,122,121,123,117,113,112,115,117,113,112,112,110,109,110,113,113,107,115,176,215,227,232,95,5,16,21,23,27,26,27,19,21,29,22,20,21,28,
147,153,136,119,89,51,67,108,133,144,142,140,139,130,108,77,46,44,53,60,60,62,66,67,69,69,72,75,81,82,82,84,90,89,88,90,89,87,88,122,80,91,93,90,92,91,103,108,102,106,111,113,120,126,136,137,154,159,163,174,175,173,177,177,177,184,187,192,190,150,87,69,83,82,83,83,82,82,77,76,72,68,72,90,107,118,120,116,115,115,115,114,118,123,117,109,110,112,116,112,112,111,111,111,111,115,115,114,111,133,205,230,150,21,14,17,21,27,27,29,20,17,24,24,18,21,25,17,
149,145,129,105,63,40,69,106,131,145,142,139,138,127,105,76,43,44,55,62,67,68,66,67,67,69,72,77,79,78,82,84,86,86,88,89,88,87,96,91,75,85,88,91,94,91,101,107,103,107,108,105,113,116,128,142,154,163,161,168,170,172,178,181,180,184,188,187,189,197,181,102,62,66,75,80,80,77,78,74,74,68,72,87,108,120,122,121,119,112,108,108,107,117,119,113,112,113,115,114,112,111,111,113,113,113,114,117,118,121,174,145,30,13,21,20,22,24,29,23,23,26,26,20,22,37,25,5,
148,138,116,83,46,44,74,105,131,145,143,140,137,126,105,74,42,43,55,62,67,70,69,64,65,69,74,75,79,80,81,84,85,85,87,88,87,95,110,77,80,78,80,88,95,96,99,100,107,109,107,108,112,117,125,134,144,150,159,167,170,176,182,182,183,186,188,187,186,189,192,188,121,81,60,72,78,77,72,74,73,66,71,87,111,122,126,125,120,113,100,96,94,106,121,117,110,115,118,114,110,112,112,113,114,116,117,118,121,131,101,26,14,18,19,26,29,25,21,17,28,27,24,25,38,31,7,63,
140,127,101,60,49,48,74,106,132,143,144,141,136,128,108,74,42,46,54,64,68,63,67,66,68,67,72,77,81,81,79,85,86,86,86,87,86,104,96,73,73,77,85,85,90,96,94,103,100,104,110,109,110,117,124,128,138,153,165,173,176,174,178,181,184,185,182,179,182,188,197,211,221,212,99,49,72,74,70,68,71,66,71,88,112,122,128,127,124,117,95,76,79,93,112,119,115,114,118,113,111,112,112,113,113,114,116,119,129,115,38,16,17,18,21,26,26,19,18,26,29,24,23,38,43,11,47,130,
132,113,78,47,50,49,75,107,129,141,145,143,139,128,105,72,45,43,56,61,65,67,66,66,68,70,73,78,79,81,83,86,86,88,87,85,90,92,74,74,78,85,86,87,92,91,92,95,97,103,106,106,106,115,113,127,137,154,171,173,173,174,178,179,173,170,181,194,203,205,209,206,212,231,189,59,56,69,68,69,67,65,70,88,109,122,126,125,124,118,100,66,52,71,100,116,117,112,114,113,112,112,112,115,114,113,117,122,125,56,15,16,17,21,27,25,24,17,23,30,22,19,30,49,35,42,112,140,
121,93,54,50,53,53,75,105,131,144,144,142,140,126,103,74,48,47,55,61,64,66,68,71,68,68,72,78,81,81,81,84,84,87,89,91,91,75,73,78,83,85,89,90,89,87,91,96,102,109,108,106,110,113,113,125,136,150,163,168,175,180,163,160,175,195,203,202,203,201,201,203,202,212,227,151,45,56,65,66,66,62,68,86,107,123,125,124,124,117,103,67,27,44,87,108,117,116,113,114,111,112,112,113,111,113,119,128,82,13,11,13,22,28,27,26,18,23,27,19,23,34,45,44,51,106,129,124,
103,68,47,55,55,51,73,106,127,141,143,141,141,127,102,73,46,46,56,62,61,66,70,68,66,70,74,75,78,83,82,87,87,86,89,91,78,73,76,80,82,87,87,86,84,87,93,99,103,111,108,109,112,116,120,123,131,143,163,164,162,149,162,189,204,202,199,196,199,199,197,200,202,205,218,225,118,38,55,64,64,61,66,85,106,124,126,125,122,120,105,75,23,21,63,94,114,118,113,113,112,113,112,112,112,115,124,103,30,27,21,20,28,27,28,23,20,32,22,20,29,43,48,57,100,130,121,117,
78,52,55,61,55,53,70,105,126,139,144,141,138,128,103,72,46,50,59,66,65,65,66,66,66,70,71,76,80,83,82,84,86,88,92,84,73,77,80,80,86,85,80,80,81,94,100,100,108,112,115,117,120,114,114,117,129,150,159,142,143,179,199,195,195,200,199,193,189,194,196,205,205,206,210,225,207,82,38,50,57,58,66,87,108,123,126,124,125,121,107,75,24,15,51,82,105,116,116,112,110,110,112,113,113,119,124,49,11,24,20,25,26,26,20,18,30,25,24,25,29,43,61,98,125,125,117,134,
57,51,57,58,55,52,70,103,125,137,142,141,137,128,103,76,47,47,59,64,67,66,65,66,67,71,71,77,80,84,81,84,86,91,92,78,81,78,79,83,85,82,86,87,90,97,99,103,109,106,112,116,115,109,111,119,132,144,124,150,183,197,194,196,193,193,188,189,195,193,194,196,197,201,203,207,217,203,122,43,45,52,61,86,107,124,125,126,124,122,109,72,25,19,31,63,92,110,117,114,109,108,113,113,118,126,81,16,10,16,26,32,27,22,15,24,27,20,27,30,34,45,94,123,127,120,135,147,
55,57,58,58,58,54,71,102,123,138,142,142,139,127,103,75,49,44,56,62,65,66,67,67,69,68,73,74,80,84,85,84,84,97,81,72,77,81,79,80,82,83,87,89,99,100,103,110,112,110,110,110,108,104,111,113,116,125,163,191,184,187,186,190,188,189,188,189,194,195,198,198,200,201,203,204,208,216,226,134,32,42,59,84,108,123,126,124,123,127,106,74,29,15,12,34,73,101,115,115,109,108,110,115,124,106,27,11,16,20,29,27,28,20,24,27,21,26,27,27,37,82,120,123,121,133,149,145,
54,59,59,60,60,56,75,105,124,136,138,140,137,127,105,75,49,44,56,62,62,65,68,65,67,66,70,75,78,82,84,78,100,110,64,70,76,82,81,78,80,81,86,93,100,103,114,113,106,114,114,109,103,103,102,102,136,162,184,190,183,181,180,179,178,187,195,194,196,197,199,198,202,199,202,198,204,209,215,218,81,26,55,81,106,120,124,124,124,120,106,77,32,17,14,14,45,85,103,112,104,103,108,117,122,54,12,18,20,24,27,28,26,20,27,23,22,27,25,25,68,124,123,111,126,144,148,146,
59,59,60,60,57,54,72,104,125,137,140,139,137,131,107,76,49,46,53,60,64,66,68,70,65,70,73,76,79,81,82,73,138,104,62,73,77,77,77,80,84,86,91,92,99,108,111,104,105,110,111,104,97,83,104,143,180,181,173,177,183,176,175,179,184,188,193,199,195,196,195,199,197,196,197,199,198,208,212,227,184,50,39,79,105,120,124,125,124,122,105,76,35,16,16,11,17,49,83,124,142,114,115,121,82,16,18,19,26,27,25,28,23,26,26,24,29,25,13,52,116,125,112,123,140,145,142,144,
61,58,58,57,56,50,69,104,124,137,139,138,139,131,105,78,49,43,54,60,59,62,67,67,67,73,74,76,77,79,71,86,168,83,68,69,75,78,78,77,83,86,93,99,105,107,110,103,107,110,100,91,84,106,156,180,172,173,176,172,164,168,182,189,189,186,189,194,196,195,194,194,193,192,200,204,200,204,207,218,235,119,28,78,106,121,122,124,124,124,106,78,35,16,18,14,0,49,160,204,200,187,196,152,28,13,21,22,28,26,29,30,28,26,21,29,25,16,37,102,128,114,118,139,142,139,138,139,
59,58,58,57,56,49,67,101,125,137,138,138,138,128,104,76,44,41,51,56,59,63,63,62,65,70,71,73,75,78,62,124,167,72,65,72,75,80,79,79,85,86,95,101,106,101,102,103,107,97,78,88,123,160,168,173,161,160,168,169,170,175,182,186,185,186,186,189,189,186,190,196,199,197,195,201,202,202,202,208,227,183,39,66,104,119,124,126,125,124,107,76,34,16,13,3,66,186,205,192,202,218,228,211,50,14,23,27,28,29,28,25,25,26,26,32,20,20,86,128,119,117,136,148,142,138,138,137,
58,58,59,60,59,52,69,100,122,139,141,140,137,129,107,72,42,39,49,59,62,64,65,64,64,67,71,70,76,76,66,161,155,73,64,72,73,82,79,83,85,93,98,95,92,91,102,105,95,80,87,135,164,164,147,154,162,159,157,165,177,175,180,181,184,184,179,176,184,191,194,196,193,194,191,194,199,199,200,201,212,226,110,53,99,122,128,128,125,124,107,72,26,7,11,101,199,186,185,211,217,216,219,238,113,9,19,26,28,26,23,24,23,24,28,25,19,63,122,125,116,132,141,139,140,140,138,137,
60,60,60,62,61,55,68,98,122,140,145,144,140,128,106,72,44,43,49,60,65,65,67,65,66,67,70,75,77,78,79,184,138,61,66,71,76,75,75,83,90,99,92,85,92,100,97,94,77,91,143,162,155,144,150,152,159,164,167,162,176,181,173,175,176,173,177,188,187,189,183,191,192,192,195,197,199,198,200,199,202,216,197,74,90,122,127,129,128,123,103,64,10,25,137,204,170,185,216,208,204,202,204,234,144,12,18,24,28,25,22,20,18,24,29,22,38,109,129,119,127,137,137,137,139,136,137,138,
61,62,63,65,63,61,70,98,123,140,145,143,142,132,109,75,47,44,53,61,64,67,67,66,66,72,71,75,79,71,91,194,129,65,66,72,67,72,82,89,91,87,88,89,102,105,97,77,94,140,150,145,144,144,148,161,166,160,168,175,169,171,175,162,160,174,181,189,186,184,186,185,192,193,185,187,189,193,196,196,199,201,214,172,105,114,125,127,126,119,87,43,73,170,199,174,193,210,206,199,192,198,209,232,145,9,22,31,25,18,18,19,22,24,17,16,80,131,122,124,140,139,137,135,137,135,133,136,
65,66,66,66,63,59,68,99,124,139,142,144,144,134,112,75,46,45,54,62,66,66,66,70,67,68,75,76,81,67,115,194,104,67,60,69,70,80,76,85,84,85,91,95,95,93,78,95,136,135,129,130,143,144,153,160,165,170,160,164,170,165,154,158,167,179,172,180,185,184,188,190,193,175,156,183,192,195,195,194,193,192,199,216,184,117,123,123,120,106,95,142,200,191,180,203,209,199,196,192,196,203,212,230,126,10,22,25,30,24,18,22,27,24,5,43,121,128,120,134,140,139,135,135,136,134,133,133,
67,67,66,67,65,63,72,100,122,136,145,147,146,136,112,77,46,45,55,61,65,67,68,66,65,66,70,75,77,60,137,178,96,74,66,70,69,67,75,81,81,91,90,88,86,80,99,133,132,122,121,123,130,152,158,160,155,154,164,167,159,152,155,171,169,169,170,171,173,181,190,191,174,159,178,184,189,190,191,191,190,188,188,193,207,148,119,115,115,148,191,196,180,188,205,203,195,195,193,195,201,207,214,226,97,11,26,22,26,23,16,21,24,18,22,93,132,122,127,140,139,138,134,135,136,134,132,131,
67,65,64,66,65,62,74,102,127,139,146,149,150,142,113,76,47,46,58,61,67,66,66,66,64,66,71,73,72,59,159,168,102,79,69,71,69,67,75,75,84,85,85,87,82,109,123,120,119,121,114,128,141,144,158,152,145,151,163,156,139,160,162,159,166,161,161,162,170,176,163,166,167,173,173,177,183,186,183,179,182,186,179,180,190,170,117,139,175,195,185,180,196,201,196,193,193,195,197,196,200,208,216,217,68,19,28,27,23,17,18,22,27,28,66,122,123,122,137,138,138,137,135,135,134,133,132,131,
66,65,66,66,66,62,75,101,127,142,148,152,151,142,115,77,47,46,57,59,63,66,65,62,62,67,67,71,66,63,183,168,112,82,68,74,71,72,77,81,83,84,91,81,101,123,123,111,115,108,118,134,141,140,135,151,161,155,140,145,159,156,160,159,156,156,164,173,175,163,160,170,178,169,178,182,181,178,173,173,176,176,174,172,172,183,170,192,187,180,191,198,200,194,193,190,194,196,196,190,197,206,220,205,38,19,23,26,24,17,20,24,31,50,106,125,120,130,140,138,137,136,135,135,133,133,132,133,
66,67,65,62,64,62,75,101,126,144,151,153,151,141,113,77,46,42,54,62,61,65,64,64,64,64,67,71,62,75,195,166,118,94,83,76,69,73,77,76,88,91,82,94,123,115,114,115,105,117,126,127,127,131,151,154,149,140,144,157,154,155,157,156,159,150,155,165,167,171,168,165,170,181,177,178,172,162,159,171,172,166,159,151,178,182,178,184,190,201,200,189,193,192,189,193,195,200,184,174,197,204,222,166,13,14,21,26,23,18,26,24,27,84,126,121,123,137,141,139,138,136,134,136,135,134,135,135,
64,65,64,64,65,62,72,101,127,144,152,152,150,142,114,81,47,45,57,62,62,66,63,64,64,64,69,70,63,79,197,161,128,107,96,81,69,69,72,82,83,73,100,112,116,114,108,98,117,126,130,111,116,132,148,146,128,149,160,146,146,156,160,153,147,151,149,152,161,159,162,171,165,175,178,163,164,168,157,160,162,147,157,180,179,171,185,195,197,197,188,189,192,191,192,194,198,192,149,152,184,191,216,104,7,19,21,28,24,18,25,21,42,117,127,120,136,140,141,137,139,137,135,136,136,136,135,136,
64,64,61,63,63,63,73,103,129,146,149,150,149,140,114,79,49,45,59,63,65,67,65,63,63,65,67,67,59,83,191,159,136,118,107,91,72,59,71,82,74,93,114,105,113,108,90,115,124,121,118,123,126,119,126,126,151,153,143,148,149,144,149,145,143,146,145,141,146,155,158,163,172,164,162,157,154,169,157,136,152,170,180,177,183,193,194,190,185,183,188,190,191,191,193,197,200,160,137,154,133,168,189,40,17,31,26,21,19,19,21,44,90,127,119,128,139,140,137,137,138,137,137,137,137,139,135,135,
66,61,63,62,61,63,73,105,130,145,149,149,149,140,117,80,48,45,57,63,66,65,63,63,64,66,67,66,54,90,190,157,135,121,107,98,70,65,71,69,97,113,100,106,102,91,110,116,118,113,114,120,129,121,121,139,135,134,149,143,143,141,138,147,137,139,140,143,147,154,153,148,159,155,153,154,146,147,146,158,171,170,176,190,199,192,185,181,182,184,189,192,193,194,196,204,183,138,154,130,127,183,146,9,14,29,27,16,23,20,30,70,123,123,121,136,141,140,138,135,137,139,137,135,136,137,135,136,
63,63,60,62,60,61,76,104,130,145,150,150,150,141,116,83,48,47,56,61,64,63,63,63,64,66,65,65,48,105,190,166,141,125,110,102,84,73,68,94,111,105,105,94,89,110,119,115,109,105,112,124,114,122,136,133,132,135,134,127,129,138,143,131,131,143,144,145,143,145,146,146,139,143,147,141,135,144,169,168,169,184,190,186,180,181,183,186,187,191,195,194,194,196,203,202,149,144,141,132,135,194,93,8,23,24,27,24,25,22,43,102,130,118,127,138,140,137,135,134,136,137,136,136,137,135,135,134,
63,63,63,63,65,65,78,103,127,146,150,150,150,141,119,83,47,42,55,62,64,63,61,65,63,64,64,63,43,112,199,176,155,136,119,116,95,62,85,106,97,106,96,89,108,112,114,108,100,101,124,112,112,135,128,112,110,119,130,117,113,96,98,142,145,139,136,137,144,142,136,137,142,138,127,134,163,169,165,177,190,188,178,176,177,183,187,189,192,196,195,195,195,199,209,177,140,131,104,84,146,196,29,12,27,26,24,36,27,24,64,125,123,122,135,138,137,135,135,134,134,135,134,135,138,136,135,135,
65,64,64,65,65,69,77,104,128,146,150,151,151,143,121,79,43,41,55,65,65,63,62,64,62,63,63,61,42,109,203,179,154,139,130,127,105,76,91,94,101,94,85,105,112,107,104,93,102,115,105,113,126,110,86,101,88,77,78,84,129,131,96,107,115,123,127,126,119,127,114,80,97,128,135,162,159,167,188,189,184,182,182,183,186,190,191,192,194,195,196,194,199,210,199,147,106,64,53,108,209,132,1,15,24,19,22,27,25,36,100,128,118,132,139,137,137,136,134,134,134,134,134,133,135,135,132,133,
66,65,66,66,67,67,80,106,128,146,152,152,151,143,119,82,46,40,52,61,63,65,65,65,64,62,62,62,42,103,201,183,171,143,111,122,112,79,86,90,90,83,103,109,105,99,91,99,104,103,106,118,114,97,110,93,80,65,45,61,137,139,111,90,78,67,82,77,62,44,38,33,30,146,156,146,169,186,189,184,185,186,183,183,188,191,192,192,195,199,196,203,202,178,124,75,50,57,92,183,195,34,12,22,23,18,23,25,19,66,123,121,122,137,141,138,138,137,134,135,134,132,133,133,131,133,133,132,
65,70,68,66,67,70,80,107,131,149,150,151,152,144,120,82,45,41,55,62,63,65,62,66,63,63,64,63,47,82,200,186,183,146,95,98,95,75,85,87,77,98,107,103,99,94,101,104,100,101,115,105,86,109,95,82,79,88,66,63,86,104,76,44,48,71,50,41,24,13,11,37,112,143,150,188,191,187,183,183,187,185,182,186,187,191,192,188,197,203,196,155,105,68,58,52,63,98,167,197,86,11,21,24,25,22,26,19,23,97,126,117,132,142,142,139,139,137,136,136,134,132,133,135,133,133,132,131,
66,70,68,61,67,70,80,106,130,150,150,151,151,144,122,81,45,44,55,62,63,65,65,66,63,64,63,60,54,57,188,195,189,150,86,100,109,91,82,76,91,107,106,97,90,96,106,98,97,111,101,88,100,97,87,90,72,57,40,31,59,89,71,67,78,57,38,56,21,5,41,131,129,152,182,186,186,182,183,180,185,183,183,184,186,188,192,197,202,168,91,56,47,52,69,85,124,180,175,54,9,18,24,20,22,26,30,17,51,121,122,125,142,143,139,139,140,138,138,136,137,135,133,133,133,132,132,132,
73,72,66,64,65,67,80,106,129,146,150,150,149,144,122,82,48,42,54,60,60,63,62,66,63,65,63,62,60,45,157,198,188,152,99,111,120,98,72,84,102,106,98,91,94,102,98,96,110,106,81,96,102,71,56,59,49,29,20,46,91,77,32,63,73,63,34,53,6,55,137,118,147,184,169,172,183,181,179,176,179,180,182,185,187,193,198,164,120,105,64,62,73,96,124,141,172,182,62,7,20,26,26,18,18,30,35,31,88,125,121,136,146,143,142,141,139,141,139,138,137,135,136,134,134,135,132,130,
72,71,70,67,65,65,80,106,129,145,150,149,149,143,122,85,47,43,52,60,62,63,64,64,65,64,63,65,64,42,111,201,181,172,129,109,115,85,78,103,105,91,83,96,97,95,88,101,101,111,91,90,56,38,55,41,28,22,23,84,80,25,41,71,58,33,21,58,71,131,118,165,185,171,166,175,173,175,175,174,178,180,182,187,198,173,111,69,76,113,118,119,137,144,146,163,179,60,5,21,29,28,24,20,20,27,22,49,115,123,121,144,145,146,146,141,142,140,139,138,136,135,134,134,136,136,131,129,
75,70,70,69,66,66,77,103,129,147,151,148,150,144,122,86,47,40,54,60,62,63,65,66,64,65,62,67,69,52,73,197,191,176,150,139,101,75,95,106,95,80,89,95,94,88,102,99,76,85,83,47,44,51,37,25,30,12,52,66,25,37,83,80,39,38,31,110,121,118,169,188,172,165,171,170,168,166,165,176,180,180,186,187,123,58,50,95,86,105,140,145,146,148,171,184,71,5,18,24,28,28,24,20,24,26,21,77,125,117,133,147,146,146,147,144,142,141,140,137,138,135,137,136,134,132,133,130,
73,74,72,68,65,66,74,101,130,147,149,148,151,145,122,86,44,40,54,59,61,60,63,62,62,61,64,69,69,67,49,143,212,173,147,156,85,88,99,94,80,94,96,88,88,97,101,96,61,45,48,48,55,37,24,60,18,24,61,27,22,46,52,51,57,61,69,119,118,175,189,180,172,168,168,170,159,164,165,178,183,179,181,127,34,50,71,91,106,95,123,138,151,178,155,52,7,15,21,25,31,30,23,19,24,23,39,99,116,117,144,148,148,146,144,144,144,143,140,139,138,137,137,136,136,133,132,130,
76,75,72,69,65,62,71,100,127,145,150,151,152,145,122,86,46,42,50,57,62,64,64,62,64,62,67,68,73,71,58,66,188,190,168,151,98,95,100,86,89,99,100,92,90,97,89,78,63,50,47,62,31,11,45,69,9,35,51,22,33,25,48,41,76,96,86,104,178,187,182,175,169,167,170,164,157,169,171,176,172,170,178,147,66,57,79,75,107,97,112,150,176,126,30,9,15,25,26,25,30,25,20,20,27,28,65,109,102,126,151,149,145,144,143,144,144,143,140,140,139,141,139,136,138,135,133,132,
76,75,70,69,66,59,66,99,127,146,151,152,153,145,123,87,44,39,50,57,61,64,61,62,63,64,66,71,73,77,71,47,125,203,185,147,99,86,80,85,99,91,85,92,94,94,87,47,42,49,65,58,26,17,51,52,28,37,21,30,42,40,48,50,69,98,109,155,172,171,176,164,163,163,162,162,161,167,171,174,173,177,185,176,106,51,68,72,75,114,120,144,92,12,14,19,19,28,29,29,30,22,18,25,23,37,87,110,103,138,152,151,145,145,144,145,142,142,142,141,141,141,139,137,136,136,132,130,
74,74,71,67,64,58,64,98,125,146,149,151,153,146,123,88,44,38,50,55,61,63,64,62,63,63,67,69,75,78,74,54,103,212,197,160,92,90,78,89,88,87,97,99,81,85,68,43,32,27,51,48,37,30,36,64,53,17,20,22,24,11,31,66,55,99,136,156,164,170,164,154,158,162,161,159,158,163,178,182,179,180,183,183,137,64,34,49,57,93,125,119,52,10,14,19,27,27,31,33,26,17,20,25,23,56,107,101,112,144,150,149,147,146,144,146,145,143,142,141,144,141,138,138,136,137,133,131,
74,71,73,69,63,57,66,97,124,144,150,153,153,145,123,88,45,40,53,60,64,64,68,65,63,64,65,71,77,81,76,56,103,213,206,113,72,88,90,84,79,100,102,95,70,34,36,46,21,18,38,50,56,34,31,50,89,30,25,17,13,20,75,73,102,134,168,168,178,173,151,144,157,170,149,148,161,176,183,186,181,183,186,185,148,75,34,20,47,76,124,124,43,17,19,19,26,30,34,33,26,19,19,21,23,84,116,104,125,138,147,147,148,146,141,142,144,143,144,143,140,140,138,139,139,136,133,129,
71,73,71,68,68,59,65,97,126,143,149,152,151,145,125,90,49,39,51,60,63,65,65,66,64,64,69,70,77,80,78,65,84,209,186,77,71,81,82,85,94,84,82,80,65,18,47,25,17,21,28,46,47,41,40,20,88,60,32,9,11,89,95,123,144,127,164,171,179,160,144,146,166,152,141,152,168,179,182,188,186,189,195,195,168,93,40,13,30,58,132,128,28,17,20,23,27,30,36,33,19,18,21,20,43,109,113,115,133,130,134,140,145,146,144,142,141,142,146,142,140,139,136,138,139,135,135,128,
70,71,71,68,67,60,64,97,126,144,149,151,153,149,124,90,50,41,49,61,65,68,69,68,66,66,62,86,97,78,79,73,64,183,169,73,85,75,81,99,93,69,55,40,35,30,55,16,27,29,22,30,36,36,59,40,61,43,6,5,82,106,125,159,141,130,154,170,172,154,154,154,140,131,146,163,173,182,184,187,188,194,197,201,184,116,49,16,15,37,113,137,40,22,23,28,29,33,38,28,18,24,26,16,68,120,109,132,139,132,130,129,130,133,136,140,140,142,143,143,142,140,138,137,136,134,133,128,
72,73,67,67,66,59,67,96,123,144,151,153,153,148,124,91,53,44,54,63,66,69,71,68,65,65,67,90,83,82,81,81,70,124,178,81,78,83,91,96,94,73,45,29,19,24,49,22,33,27,25,26,29,26,68,63,59,71,0,68,108,124,163,163,153,136,152,182,172,152,149,130,126,142,151,169,176,182,187,189,189,196,198,200,191,138,59,21,9,26,94,143,51,26,26,27,33,35,39,23,19,26,22,25,96,118,115,143,145,137,134,131,129,127,131,129,129,134,135,141,141,138,136,135,135,133,130,126,
72,72,66,65,63,55,64,95,123,144,152,154,154,147,125,91,52,46,59,62,66,67,68,67,68,68,69,81,81,81,86,85,78,85,154,91,79,98,98,100,71,34,27,52,19,16,47,33,34,28,22,29,37,23,47,37,29,73,53,106,110,150,159,177,169,125,157,182,153,140,130,129,143,148,153,165,178,179,185,191,190,195,198,200,201,155,74,30,15,18,76,145,54,18,27,32,32,35,34,25,22,27,18,51,118,114,127,149,147,145,142,139,136,133,133,130,126,126,127,129,130,132,132,131,132,134,130,126,
69,69,67,65,64,58,61,96,123,145,153,156,155,147,126,89,49,45,55,62,67,66,71,71,67,67,72,77,82,80,80,79,82,88,88,83,90,103,101,89,37,33,21,51,29,20,21,47,51,18,18,35,36,29,31,52,0,49,104,105,143,137,153,175,175,141,166,162,135,133,131,138,147,150,154,161,174,182,183,184,188,192,196,201,200,174,91,45,17,16,57,143,65,20,27,32,36,39,28,22,26,22,21,85,119,111,137,148,143,143,143,148,145,146,138,136,131,127,128,126,122,122,123,126,130,133,130,129,
68,68,66,63,63,57,62,96,126,145,151,155,156,149,126,86,50,42,53,62,67,68,68,68,68,66,72,76,81,83,83,83,100,99,95,112,85,100,94,66,36,50,17,69,22,20,43,60,30,15,22,37,29,47,39,35,20,81,89,147,152,141,148,178,177,174,146,110,122,136,142,147,153,155,154,157,168,178,180,180,184,189,193,198,200,185,104,37,14,15,39,139,83,28,37,33,37,38,26,25,27,20,40,105,112,116,141,146,144,143,142,145,147,150,145,139,137,133,130,127,125,123,122,122,121,123,123,127,
67,67,66,65,64,58,62,95,124,143,152,155,156,148,127,90,51,45,53,61,66,69,69,67,66,68,70,77,81,85,79,127,129,41,14,81,138,87,66,32,62,33,34,76,13,24,34,29,18,20,28,35,34,47,37,14,73,91,139,160,169,141,145,185,190,136,70,66,75,79,97,130,155,161,155,151,160,174,180,173,178,185,190,200,189,149,77,20,12,12,33,128,101,27,37,34,42,35,22,24,27,20,63,116,108,127,144,141,140,140,140,140,143,144,144,139,136,137,136,133,129,129,127,122,120,121,118,115,
69,68,69,67,65,59,61,93,124,144,152,154,157,150,128,91,49,46,56,61,66,71,67,67,66,67,70,76,80,84,94,125,98,13,9,96,118,60,37,41,61,20,60,75,13,29,39,42,33,19,15,42,61,44,16,45,104,124,158,172,174,133,172,187,130,99,114,115,103,64,40,47,85,137,152,147,153,170,175,171,175,179,172,136,97,72,62,40,16,15,24,113,121,28,37,40,37,29,24,24,29,23,82,115,109,134,144,140,137,138,137,136,138,139,141,138,135,136,138,136,136,136,132,126,125,120,116,111,
67,70,72,69,65,56,59,93,123,144,153,153,157,152,129,93,50,46,54,63,68,68,66,65,63,66,68,69,72,97,127,115,121,90,67,88,71,38,30,66,41,54,42,57,29,36,22,37,58,10,12,20,48,30,17,93,122,159,163,187,157,158,181,106,73,87,87,79,107,77,72,59,52,84,128,136,144,166,177,172,172,152,100,67,61,69,72,52,31,16,23,104,125,37,33,38,38,24,24,28,25,37,102,110,116,141,139,137,136,136,137,134,134,138,139,137,135,133,135,136,138,138,135,132,132,124,118,112,
67,70,69,65,63,53,56,94,124,144,154,156,156,150,130,95,52,41,51,59,66,67,65,64,63,62,59,87,121,117,127,126,132,120,98,28,26,47,64,73,43,75,28,36,38,42,20,14,66,45,15,16,13,9,68,109,155,158,181,187,172,167,75,34,38,30,24,21,26,13,44,87,90,86,106,123,136,166,180,183,169,99,57,34,20,24,30,33,28,13,24,98,128,48,31,39,30,21,23,27,16,53,117,108,126,141,138,135,134,135,135,133,135,135,138,135,133,135,133,134,136,136,132,127,128,124,120,116,
65,64,63,60,59,49,49,88,122,145,155,156,156,148,126,93,50,39,50,57,61,67,62,61,60,49,79,172,147,106,123,120,105,50,32,10,62,58,64,51,61,88,29,31,29,59,29,11,25,78,47,18,7,32,102,140,159,163,189,188,171,70,18,18,17,17,11,42,102,44,4,44,97,92,100,114,131,169,195,190,89,22,23,53,57,17,25,26,19,15,22,90,131,52,37,40,24,21,25,27,17,74,119,115,138,139,136,134,132,132,131,135,132,135,134,134,134,134,133,131,133,132,126,124,121,119,119,114,
65,63,61,59,54,45,45,89,123,149,157,156,159,152,126,91,47,42,53,61,65,63,65,65,59,45,84,171,130,110,125,101,85,26,20,54,45,43,29,36,86,73,24,21,15,46,56,14,16,25,32,28,14,75,117,160,158,176,197,185,90,36,17,24,49,35,29,55,182,168,57,48,75,83,94,107,131,176,211,131,24,24,35,92,128,37,16,22,20,19,25,83,133,56,48,38,23,23,26,20,33,100,119,122,140,137,136,133,130,132,131,131,132,130,131,133,131,132,130,129,129,126,122,119,114,112,110,113,
67,64,63,62,56,46,44,87,122,147,157,160,162,153,126,92,54,45,55,66,68,67,68,73,66,29,43,109,147,195,126,44,22,12,53,47,31,43,36,60,87,83,20,21,20,27,54,19,18,21,13,10,47,84,135,147,168,193,189,109,77,78,49,25,77,62,45,106,202,196,109,68,72,79,88,105,138,191,199,86,72,60,51,106,141,48,13,16,18,18,30,81,139,59,56,33,24,26,26,18,48,116,115,129,139,136,134,132,132,130,130,130,132,132,131,132,129,127,128,126,126,120,117,112,108,112,124,142,
69,66,66,61,58,44,44,86,122,146,158,160,160,155,130,91,55,50,59,68,73,73,75,38,29,66,100,145,181,166,60,31,21,63,71,25,35,54,54,81,83,98,38,25,17,17,26,26,21,23,9,22,85,122,154,166,195,186,105,77,90,109,101,64,69,90,106,160,179,165,123,94,87,81,89,99,140,205,189,85,95,96,112,152,106,33,26,22,23,28,36,70,145,67,56,29,21,23,28,20,70,118,116,135,137,135,133,130,128,132,140,132,132,135,131,128,129,125,124,121,119,118,110,114,131,147,161,174,
70,71,68,59,52,43,42,86,124,145,157,163,165,159,133,95,55,49,61,69,77,77,87,30,77,131,116,122,105,27,16,69,79,69,52,11,47,58,48,71,102,100,76,29,16,20,19,19,24,16,4,60,95,152,159,185,191,97,69,98,103,108,113,108,96,80,86,104,100,127,140,116,86,89,88,96,133,200,198,138,112,103,98,84,41,40,46,24,19,30,37,61,151,80,50,25,21,22,26,40,99,112,122,140,137,132,131,131,128,130,136,132,130,131,132,126,123,121,118,116,111,115,129,150,168,176,179,177,
68,69,64,57,50,42,37,82,122,146,158,162,164,159,133,98,54,45,60,68,74,69,88,117,127,111,58,54,49,19,20,31,96,106,80,27,34,50,69,60,82,107,78,28,19,21,19,23,22,8,28,98,115,156,173,196,100,53,87,104,115,120,117,118,112,106,102,110,118,130,129,119,91,97,90,88,127,193,205,154,122,103,95,83,62,70,55,25,14,26,34,57,155,88,41,25,20,30,20,44,114,109,129,139,134,133,130,130,132,130,127,130,130,130,127,124,121,121,115,111,117,144,169,180,181,179,178,178,
66,59,58,49,49,33,30,79,121,143,156,163,165,159,134,98,55,46,58,68,74,70,76,106,100,70,59,63,31,24,47,62,73,67,62,14,28,54,52,99,72,78,77,23,18,19,17,24,25,15,78,92,147,173,200,115,42,75,90,105,119,126,135,135,135,132,133,143,144,142,141,118,101,102,89,88,122,187,208,171,142,125,107,94,85,81,64,28,19,30,31,50,155,94,35,26,20,24,16,64,115,112,135,136,134,130,129,130,131,131,129,128,128,128,125,122,121,119,109,118,155,182,187,185,181,179,178,178,
60,61,53,50,45,30,32,77,120,144,157,159,163,157,133,98,55,46,58,63,72,87,99,105,120,102,97,48,27,43,69,88,77,76,32,11,27,66,68,81,92,106,74,50,28,23,20,23,18,45,96,112,171,196,140,27,60,82,90,102,117,125,138,143,151,149,149,149,147,151,136,115,108,101,92,84,112,181,210,173,150,128,109,100,91,84,70,29,21,32,28,38,153,106,25,22,22,23,21,87,113,121,140,136,133,131,131,131,131,132,129,128,126,124,123,119,118,112,119,156,183,190,188,183,180,178,180,181,
56,58,49,48,42,30,31,79,120,146,155,158,163,157,134,97,54,43,54,73,93,105,112,106,71,47,46,30,39,58,70,94,98,48,21,19,16,27,57,76,62,20,84,98,35,20,22,20,16,86,95,147,190,175,30,32,73,84,90,100,113,122,137,147,153,154,154,154,154,149,135,120,113,104,93,87,106,173,214,176,142,132,111,97,91,90,71,28,24,38,31,31,142,118,26,15,22,19,31,106,113,127,141,136,133,133,132,130,129,130,128,125,126,124,123,118,112,113,149,180,186,187,186,184,181,180,185,188,
50,48,42,44,43,31,29,77,119,145,155,159,160,155,132,96,55,46,57,73,77,81,79,57,64,62,49,35,71,46,85,99,53,33,20,24,24,24,33,36,30,11,81,113,50,12,17,11,40,100,118,181,189,71,8,48,78,85,89,96,109,119,128,144,152,157,159,151,151,144,130,117,112,107,94,89,105,166,217,181,140,130,118,100,92,92,64,26,22,33,35,25,132,126,31,15,30,14,51,113,117,138,141,132,136,133,129,129,128,126,126,127,124,124,121,115,107,133,176,188,183,184,184,184,185,189,194,196,
47,43,44,40,37,28,28,74,119,141,153,155,156,152,131,100,52,45,64,67,68,77,76,97,80,66,66,73,51,27,65,93,52,29,24,28,25,21,30,35,24,20,71,97,111,27,10,8,76,91,157,204,126,13,25,45,76,84,92,97,105,115,122,132,143,153,157,150,146,138,125,108,106,103,87,90,104,149,212,185,138,129,119,105,95,88,56,22,20,35,31,16,130,134,50,12,33,22,73,115,124,150,137,135,133,133,129,127,125,126,126,124,123,122,118,109,116,163,186,184,181,183,185,188,193,198,198,196,
47,44,47,44,37,25,27,76,119,140,152,152,155,151,128,98,51,41,86,68,86,114,101,45,65,97,72,40,50,52,75,109,72,31,35,27,17,16,31,51,26,32,108,82,93,83,3,29,95,107,198,179,28,17,29,41,70,83,91,95,103,114,123,129,137,147,147,146,142,135,123,103,98,97,87,84,98,142,206,194,137,126,115,102,95,87,44,17,27,39,34,12,117,133,68,14,24,25,97,116,130,144,138,135,135,131,129,128,127,126,124,123,121,120,115,109,143,182,187,183,181,184,189,197,203,202,195,193,
48,48,46,44,34,23,23,73,118,140,151,151,155,151,131,97,49,36,76,96,104,100,65,36,93,75,59,39,73,76,91,104,88,38,31,24,11,18,45,68,36,69,130,128,34,48,0,66,95,152,202,68,0,24,39,39,67,84,90,93,100,110,119,125,129,134,139,141,139,134,119,101,94,90,85,81,94,134,196,209,137,125,114,104,95,80,32,17,29,45,33,8,103,143,75,13,17,42,111,115,136,141,134,131,134,133,132,129,127,128,125,123,118,119,109,120,169,188,184,181,183,190,198,202,203,201,197,195,
48,47,45,44,33,19,17,71,116,141,152,153,156,153,134,97,51,36,55,85,84,99,66,46,66,69,56,53,78,61,70,113,73,37,17,27,20,18,48,50,89,84,62,71,17,10,29,84,104,184,112,3,10,30,50,39,65,81,89,94,97,106,115,119,123,125,133,136,133,125,110,91,85,97,88,83,94,125,186,218,140,119,115,101,94,71,22,19,30,43,32,5,90,142,94,18,12,66,119,119,137,138,134,131,131,130,131,130,128,128,125,124,120,114,109,146,185,187,184,183,189,199,203,200,198,200,201,199,
53,49,47,41,31,18,16,70,116,143,152,154,157,156,134,97,51,51,87,81,75,83,47,48,73,77,49,47,77,39,76,105,72,53,24,32,24,15,47,73,58,88,47,16,7,31,126,113,120,156,56,6,12,34,57,39,67,82,89,92,97,105,110,117,120,125,127,131,132,121,110,76,86,105,108,95,87,120,182,213,134,113,110,96,91,52,15,21,29,46,31,5,70,147,109,23,12,90,123,124,141,135,133,130,130,129,128,129,128,128,126,125,118,108,119,169,191,185,184,185,195,202,201,197,198,201,201,200,
54,49,48,41,34,23,25,77,117,142,150,152,156,155,134,98,64,59,64,63,75,81,45,51,92,73,23,77,69,34,71,99,94,73,33,28,37,12,28,31,45,72,18,11,0,83,173,169,170,90,8,12,14,32,60,44,67,82,87,90,96,104,109,116,118,120,125,128,129,123,110,84,93,76,59,77,76,99,161,180,125,114,109,98,80,24,17,25,32,40,27,8,54,146,111,31,23,106,123,131,139,134,132,130,129,128,130,127,127,126,125,122,117,108,135,179,188,184,185,193,198,199,199,201,201,203,204,200,
48,46,44,42,35,32,42,90,122,141,150,152,156,155,135,101,55,40,55,64,77,72,52,54,77,49,34,95,55,49,71,92,112,84,34,20,52,45,8,19,90,45,19,25,27,106,150,179,114,6,17,20,14,33,70,51,70,80,85,91,95,103,111,114,116,118,124,126,130,126,118,96,85,74,66,67,67,84,145,157,125,112,104,98,54,19,23,25,36,42,31,13,36,140,118,39,48,120,123,134,138,134,131,128,129,131,128,128,125,124,123,121,114,111,149,184,187,186,192,199,200,200,201,204,204,204,202,200,
47,46,45,42,37,40,56,99,127,142,147,147,155,158,136,101,55,42,58,64,79,79,30,50,45,28,77,53,52,55,80,80,105,112,54,4,65,116,12,30,56,33,59,96,117,77,116,154,23,10,40,29,13,38,78,52,73,81,85,89,92,98,107,110,112,115,121,125,129,127,123,115,101,91,100,104,107,159,174,145,124,112,102,89,31,21,24,28,46,51,32,18,22,129,121,46,68,125,125,138,136,134,131,130,127,129,129,127,126,126,123,120,113,117,162,188,186,188,197,202,200,199,202,204,204,204,201,202,
48,44,46,43,35,37,66,106,130,141,146,150,155,156,138,102,58,44,56,61,84,102,32,41,49,85,56,22,46,59,80,87,81,115,94,29,52,81,32,27,40,99,117,159,94,76,163,68,17,29,31,34,18,38,81,57,75,84,87,89,94,101,104,107,108,116,122,124,128,128,123,120,115,108,124,163,147,184,179,144,118,109,103,65,22,23,25,34,49,49,36,27,16,117,120,55,93,124,126,138,135,134,130,130,129,127,127,126,126,126,123,120,111,123,171,187,186,193,201,201,199,199,202,203,204,205,203,205,
44,41,40,39,31,34,69,105,129,142,145,147,156,156,138,104,58,41,50,67,103,85,36,51,91,50,35,28,43,46,51,78,62,100,110,60,73,39,19,28,90,136,172,138,52,114,93,8,24,21,28,37,19,27,78,65,73,82,87,89,93,101,104,103,105,110,115,118,118,125,119,118,118,120,149,192,160,185,181,140,114,109,96,33,22,23,25,38,49,44,33,23,9,101,123,71,108,121,130,136,134,131,128,129,128,128,124,126,125,126,123,119,109,130,177,186,190,200,203,200,200,200,200,203,205,205,205,205,
41,38,36,36,32,39,63,102,127,140,148,151,157,159,141,105,56,38,53,93,84,78,38,74,72,20,45,45,44,50,42,63,48,78,108,106,62,9,56,77,91,152,167,73,82,109,15,28,28,20,25,42,21,20,73,64,66,81,87,90,92,99,104,103,102,101,108,113,113,117,114,114,123,129,157,197,173,187,183,137,105,111,72,17,25,26,28,39,50,42,34,25,10,90,121,82,113,120,134,135,134,132,129,127,127,129,126,124,125,124,121,115,107,135,181,189,196,203,201,200,202,201,201,205,207,206,205,205,
35,29,35,37,30,37,59,102,131,143,148,151,159,160,141,105,54,33,81,81,69,79,26,61,63,30,39,40,55,68,58,51,61,45,77,118,54,39,99,154,168,177,91,65,124,34,12,50,25,19,28,46,25,18,66,59,58,78,87,91,91,98,102,105,101,103,100,95,105,107,111,108,114,115,114,130,150,127,127,105,98,105,38,17,30,25,29,41,49,46,39,26,3,80,122,93,117,121,135,135,133,130,128,127,130,128,129,124,125,122,120,115,104,138,181,194,202,204,201,202,202,202,203,206,208,207,206,206,
28,28,34,34,29,36,63,106,132,147,153,155,158,158,140,101,48,63,88,53,101,80,26,41,41,40,43,29,54,99,81,65,51,71,75,71,67,102,114,183,208,114,56,124,75,9,18,33,21,19,28,41,29,18,60,53,51,75,88,92,87,93,99,106,109,111,75,58,64,74,78,77,68,60,59,73,81,58,71,78,112,80,18,22,25,23,34,40,45,49,30,34,9,65,120,109,121,123,135,137,132,132,129,128,128,128,128,126,124,123,122,113,105,145,185,200,204,203,203,201,201,203,204,206,209,209,207,208,
27,29,31,31,30,46,73,107,131,148,155,155,161,158,137,95,77,96,49,70,111,69,39,33,23,36,45,39,60,117,68,79,74,70,77,51,66,110,96,188,170,63,107,122,19,23,19,27,25,21,30,35,35,22,53,53,50,70,84,87,86,91,96,101,113,111,96,82,70,67,71,83,88,99,105,124,133,96,98,111,107,36,18,25,22,25,33,36,49,47,30,43,16,49,128,120,121,127,137,136,132,133,133,130,127,125,129,126,125,125,121,112,106,152,192,206,207,205,204,203,205,205,205,208,208,208,207,206,
28,29,30,31,27,50,69,105,131,144,155,159,163,157,142,113,97,49,43,100,84,58,50,66,16,27,52,45,74,127,42,64,84,69,45,76,114,114,94,160,93,111,141,40,22,29,20,21,26,20,30,33,36,25,42,50,44,65,76,81,82,87,90,98,108,112,111,98,88,85,82,85,105,133,141,143,144,105,114,120,66,14,21,25,18,24,26,33,54,49,31,46,20,46,133,126,125,128,138,138,136,134,133,133,131,130,128,125,127,124,120,110,105,158,201,209,206,204,206,206,205,207,209,209,206,204,203,201,
27,24,25,27,25,48,66,99,129,144,157,160,162,158,144,116,54,28,81,97,73,41,71,67,14,43,54,47,101,112,72,65,59,86,90,91,122,115,111,150,113,161,55,22,30,32,30,26,27,26,32,36,41,27,46,49,39,56,71,74,79,84,92,95,101,106,108,103,95,88,88,82,85,93,96,88,94,113,120,96,29,19,24,25,24,27,24,37,51,50,36,46,24,45,133,129,129,132,139,136,135,136,134,133,131,131,128,126,126,122,120,109,104,164,208,210,207,206,207,209,209,210,208,202,199,198,197,197,
26,23,24,22,27,58,61,93,121,141,157,159,161,159,138,100,50,34,100,75,70,27,82,54,14,52,39,35,129,99,87,105,56,70,117,89,86,98,125,159,162,77,20,30,28,32,26,27,25,31,33,32,36,26,38,48,37,43,61,67,73,80,87,94,95,102,106,102,98,94,92,91,86,85,87,95,117,115,109,49,20,19,21,28,34,27,22,43,52,55,36,44,29,42,134,131,127,133,138,136,135,135,135,137,135,132,130,127,126,123,119,105,100,167,212,213,208,208,209,210,210,206,202,199,201,203,203,202,
26,23,21,17,35,74,70,94,116,138,156,157,159,158,140,105,52,33,89,74,53,40,65,34,19,50,35,32,127,110,90,119,91,74,86,84,69,90,138,195,105,16,27,24,27,30,26,26,27,26,28,31,33,31,25,39,36,39,48,63,70,77,86,91,97,102,102,104,103,103,105,116,123,127,122,126,123,114,77,26,24,20,26,31,34,26,19,46,54,53,40,47,31,37,133,139,125,137,139,137,135,136,134,134,135,132,131,127,124,122,117,103,99,170,214,216,210,210,210,209,207,204,204,205,205,203,203,204,
21,22,22,21,45,73,73,95,116,138,154,156,157,156,138,103,54,34,70,79,50,57,58,26,20,53,27,36,94,84,88,112,104,78,63,92,83,70,121,149,27,22,28,28,26,34,22,27,26,24,20,28,30,28,24,34,31,33,31,43,61,68,80,91,98,100,104,108,110,124,126,126,143,145,137,132,121,121,42,23,22,23,29,36,32,29,20,55,59,56,41,48,34,33,136,140,127,139,140,138,135,135,132,133,136,132,130,126,123,122,115,103,103,181,216,215,210,207,206,206,208,207,207,205,202,200,202,200,
21,24,20,22,44,69,69,96,116,141,155,156,158,157,140,103,53,35,64,67,36,45,68,29,28,47,25,38,96,64,35,85,116,106,86,100,102,68,81,73,36,27,28,24,31,34,22,30,25,27,21,22,30,29,28,31,33,36,33,17,34,53,67,88,92,99,103,113,116,127,142,139,142,141,146,139,124,101,20,30,29,29,30,36,25,29,21,58,63,56,45,45,37,35,135,140,127,138,141,136,132,133,133,132,133,132,130,125,122,120,114,102,110,193,218,212,206,205,207,209,209,205,202,199,199,200,199,187,
22,24,20,20,34,58,77,99,118,141,153,155,158,158,141,104,52,28,66,51,22,46,66,32,37,42,25,24,106,88,32,62,90,107,120,103,122,91,68,42,30,28,28,26,31,37,24,33,26,30,26,21,26,30,31,30,34,34,42,25,16,26,47,64,73,87,94,103,112,117,130,139,143,137,138,130,117,80,19,32,35,35,33,39,29,24,25,62,65,54,50,50,44,37,134,139,124,127,132,131,132,133,134,132,131,131,126,124,121,119,114,96,124,203,219,210,204,207,210,209,206,201,199,200,191,164,122,78,
19,21,19,18,25,56,72,92,121,142,151,152,156,156,138,99,41,75,107,76,25,50,44,34,39,32,25,17,97,122,62,47,80,92,90,102,136,117,124,103,24,23,28,28,38,44,22,34,27,24,28,24,21,27,34,34,37,31,41,43,29,32,41,47,60,72,83,90,100,112,121,130,139,130,126,116,111,68,18,26,35,34,34,37,30,24,29,62,68,58,55,54,43,47,137,132,103,96,108,114,120,124,129,130,131,129,126,124,121,118,110,94,143,209,215,207,204,205,206,204,201,196,186,153,101,44,14,12,
24,26,16,15,21,48,55,87,120,139,153,153,152,155,134,87,102,147,66,80,27,40,46,37,38,32,23,18,83,124,97,41,45,77,98,92,119,119,65,120,114,27,20,25,39,44,19,35,24,24,26,23,23,23,34,32,31,25,29,47,54,72,86,94,99,106,103,107,109,121,131,128,133,136,139,147,161,149,106,61,31,28,27,33,25,26,30,60,67,62,52,55,41,54,138,118,86,84,85,93,99,102,107,113,121,125,124,123,121,113,105,97,165,213,208,201,204,203,200,200,194,175,134,55,11,13,23,35,
36,34,25,19,20,39,43,81,114,138,150,149,151,150,129,133,132,52,49,68,12,35,55,34,34,50,44,23,63,106,109,73,41,98,127,70,82,110,66,69,143,108,28,24,43,43,20,41,28,25,24,26,22,27,27,32,30,26,25,49,66,87,96,92,96,99,102,107,108,116,120,116,115,117,132,155,176,192,197,181,131,70,28,21,24,24,34,65,66,58,52,55,45,64,137,109,95,99,89,87,85,84,85,89,94,100,105,108,113,109,100,100,175,210,201,197,201,202,202,192,180,148,68,15,18,31,46,54,
87,62,40,28,27,30,26,58,103,136,148,148,148,154,155,135,48,45,99,43,11,21,46,40,20,44,65,41,28,70,100,80,84,125,85,61,77,95,76,112,112,90,83,17,37,37,22,42,27,23,22,28,23,23,26,35,32,29,24,45,71,86,89,90,90,96,103,102,106,109,109,109,111,117,137,159,177,185,188,194,199,190,138,61,12,10,27,61,64,53,47,51,36,67,137,111,110,113,109,100,95,88,81,76,74,75,81,82,83,88,81,84,170,204,196,197,200,201,202,188,141,57,18,23,34,47,56,58,
119,109,79,51,44,31,20,48,97,136,145,148,148,157,147,99,58,108,93,10,18,16,40,71,7,32,83,62,38,17,90,89,77,94,55,87,84,97,104,106,111,45,93,49,30,34,18,42,27,24,21,29,32,24,27,31,39,34,23,42,69,82,86,89,92,93,101,101,105,106,107,110,116,124,145,165,176,179,183,186,191,194,206,192,109,19,18,53,60,50,45,45,34,70,132,116,123,119,119,111,111,106,99,89,83,72,70,65,74,93,70,55,161,203,196,202,200,199,188,145,57,16,40,46,49,55,57,56,
120,127,120,90,67,43,15,47,98,134,147,146,149,151,136,103,122,99,44,16,16,10,57,89,56,79,70,53,37,51,52,65,96,52,46,71,98,107,128,104,71,78,51,93,33,28,25,46,30,28,24,30,38,30,26,32,41,42,25,42,71,81,82,90,91,95,102,109,109,105,102,109,120,134,146,161,172,174,178,180,187,191,195,203,210,143,30,30,54,42,43,48,25,80,130,122,129,123,122,119,118,115,111,105,98,91,85,72,83,106,72,63,172,206,201,207,203,198,137,42,18,49,53,49,59,66,59,54,
115,131,139,125,93,54,20,43,98,139,153,150,151,154,131,132,163,71,31,21,21,21,35,37,68,58,33,39,61,64,23,89,45,38,49,72,76,110,123,136,51,89,84,92,52,20,25,43,30,29,28,31,38,29,30,41,42,60,26,34,71,83,89,86,90,105,101,105,108,104,105,114,126,135,142,153,162,166,172,178,182,186,193,197,202,215,150,35,37,33,43,46,23,86,129,123,130,126,124,124,122,118,116,114,108,105,100,90,95,106,76,100,193,207,206,205,202,181,84,11,48,64,55,56,73,70,59,60,
92,118,139,141,127,78,20,43,99,138,155,156,154,155,130,138,133,81,21,21,28,29,44,29,33,27,46,37,23,33,25,72,52,38,48,66,74,88,126,114,99,77,120,75,87,17,27,44,34,29,28,31,40,31,31,41,48,75,37,25,73,86,82,89,98,103,104,106,107,106,111,119,128,136,140,147,155,159,165,170,178,184,189,195,199,205,219,135,23,19,37,42,25,96,126,124,130,127,123,122,122,120,119,116,113,109,107,102,102,108,89,136,203,207,206,206,193,144,51,36,63,60,60,72,84,69,59,68,
39,94,134,155,147,99,25,40,101,141,156,156,158,157,134,131,115,40,17,18,19,35,38,31,19,27,70,42,21,36,47,28,69,42,48,49,70,89,105,110,132,92,64,99,110,21,17,38,32,25,22,26,39,29,21,32,50,86,48,21,67,77,91,98,96,103,106,105,104,107,111,117,123,132,136,143,153,155,160,167,175,181,187,192,197,203,209,217,94,8,28,29,22,105,120,125,128,127,124,124,122,123,120,117,115,112,107,106,108,112,101,161,210,207,207,206,182,95,41,60,63,63,71,84,75,63,66,75,
12,58,130,160,154,117,31,31,102,139,156,156,158,156,138,115,119,56,16,19,23,46,24,30,22,35,77,37,29,15,50,39,51,56,63,74,56,75,87,104,142,107,15,81,146,32,12,37,36,25,22,27,42,31,24,25,56,87,51,17,61,83,94,98,97,98,104,107,107,108,110,117,121,129,136,140,146,153,160,166,175,179,185,191,194,198,206,220,191,33,19,21,22,112,117,127,126,124,124,124,120,120,118,117,116,113,109,102,102,119,137,182,210,209,206,204,160,59,48,61,65,72,81,75,57,64,74,75,
8,33,119,165,159,125,28,26,101,139,158,157,157,158,142,105,98,59,16,20,32,32,22,26,18,44,84,28,40,12,25,55,53,41,62,85,79,56,79,129,138,78,17,84,172,32,14,36,44,29,21,27,35,23,25,30,67,75,51,23,61,85,93,91,98,99,103,106,107,110,115,116,119,126,132,136,144,151,158,164,172,177,184,191,196,201,203,210,223,109,4,9,23,122,119,131,127,125,124,122,120,118,115,116,115,112,104,97,117,159,183,198,210,209,207,194,118,54,61,63,69,81,79,63,58,70,73,75,
8,31,110,159,163,121,25,26,100,140,160,159,159,161,144,116,110,57,18,25,33,26,21,26,16,71,87,17,38,25,30,32,27,37,57,80,78,55,70,125,127,104,16,77,145,17,18,45,45,30,25,26,36,21,22,40,67,77,64,22,64,86,96,93,99,104,102,101,104,107,113,113,119,124,127,133,143,148,156,163,170,175,183,191,195,200,203,207,220,182,21,2,33,123,124,130,130,128,126,122,121,119,113,113,113,106,99,108,166,192,192,204,212,209,204,168,78,57,62,68,78,84,70,60,67,72,73,78,
5,17,100,155,163,126,27,22,99,142,159,159,160,161,142,118,105,28,24,32,21,18,19,15,25,104,74,18,24,34,30,24,24,27,43,69,91,37,67,126,127,104,71,106,134,72,15,42,38,29,27,23,28,30,27,52,79,90,67,26,67,89,95,99,101,99,100,101,101,105,111,113,115,121,127,133,139,144,153,159,169,174,181,189,196,200,203,206,212,220,74,0,48,119,128,129,126,125,125,122,119,118,114,112,107,107,95,137,206,208,198,206,212,211,194,124,61,58,59,71,81,81,63,58,73,77,76,74,
6,15,90,157,166,131,34,18,96,143,158,158,161,161,144,117,80,26,34,20,20,19,18,23,68,76,54,17,26,42,23,14,30,26,36,45,94,65,87,126,119,104,120,142,74,42,27,29,31,30,31,28,24,26,39,73,91,91,57,34,70,88,94,101,103,104,101,101,103,105,108,112,115,119,127,132,135,141,151,158,165,176,182,186,194,197,201,204,206,224,130,0,57,119,130,128,126,125,124,121,120,119,115,113,108,102,93,159,212,210,201,209,212,207,168,93,66,63,61,75,84,70,61,68,77,76,72,64,
5,12,88,155,165,136,46,18,93,140,156,155,155,154,141,116,91,40,23,21,22,22,32,46,28,50,62,24,30,39,22,20,32,27,49,34,36,94,117,120,88,71,114,130,86,70,58,40,37,40,28,29,21,27,48,81,91,91,52,35,74,90,97,96,104,107,103,102,100,103,107,109,112,117,123,130,134,138,146,153,163,174,181,186,193,195,199,203,206,215,180,10,61,122,128,129,124,124,121,119,120,120,116,112,107,102,102,171,212,201,200,210,211,195,133,86,72,65,67,77,82,66,62,72,76,73,64,58,
6,9,77,151,166,142,50,18,91,139,156,156,156,159,142,119,95,34,21,22,22,24,28,31,24,44,52,27,32,29,30,20,28,33,60,25,19,74,110,106,101,51,25,44,48,55,72,81,86,59,28,26,22,36,59,85,92,93,49,45,81,93,98,99,105,105,104,102,97,101,104,109,110,118,122,128,132,135,144,149,162,170,178,185,190,193,196,201,204,208,206,51,66,123,128,131,124,124,121,120,119,121,118,113,106,103,108,177,211,199,199,212,209,172,100,82,75,64,68,75,72,57,62,78,72,66,63,66,
9,10,65,146,165,146,55,23,90,138,156,159,159,160,145,124,90,24,25,20,19,22,29,39,25,36,40,32,23,32,34,15,26,33,61,38,55,68,90,96,89,110,48,40,12,22,30,35,39,53,35,19,25,48,69,88,95,92,39,58,88,97,100,103,105,105,107,102,99,101,104,106,110,114,118,126,130,136,144,148,155,167,177,183,189,192,196,199,203,204,216,100,69,125,132,129,123,124,121,121,121,119,119,113,109,107,107,158,200,192,199,214,204,149,85,80,75,64,65,68,52,59,72,75,69,68,65,71,
15,8,53,137,164,146,68,27,87,136,155,157,158,157,142,124,104,39,26,17,23,42,49,28,22,37,35,29,32,30,37,24,31,46,43,58,41,95,107,104,51,82,105,76,42,24,27,28,29,24,28,18,34,56,75,89,95,79,35,66,92,99,105,106,108,107,104,103,102,102,103,104,109,113,118,123,127,134,140,144,152,163,174,180,186,190,196,198,202,203,213,154,87,121,118,124,125,125,127,126,124,122,119,115,112,113,112,119,148,169,204,213,198,133,78,72,65,62,67,56,46,74,74,67,64,68,71,67,
14,8,45,133,160,147,82,30,85,135,154,156,158,159,143,121,109,49,29,18,34,40,27,21,26,40,35,34,39,33,34,25,38,48,18,69,48,42,59,100,55,39,105,144,52,19,22,29,24,21,19,19,41,66,82,90,93,56,38,79,96,103,104,106,109,108,104,106,105,101,101,105,109,113,118,121,124,129,134,140,151,161,169,176,185,189,194,199,202,203,205,193,115,99,83,95,105,115,122,127,128,127,126,119,118,124,121,114,107,154,212,214,185,111,75,70,57,64,62,47,60,77,70,62,63,71,71,51,
11,8,42,128,161,152,83,32,81,133,153,156,158,159,144,115,92,55,30,17,27,24,22,26,36,37,32,49,35,20,28,15,35,33,31,79,94,33,17,52,54,49,81,90,19,25,20,25,20,14,21,33,50,75,82,90,86,36,50,92,100,102,105,107,109,110,107,107,105,102,103,104,108,114,117,121,124,127,134,141,148,153,164,176,182,188,194,200,202,203,206,212,135,53,52,56,68,80,91,104,113,115,120,124,127,136,121,106,113,173,215,210,163,92,66,53,57,66,45,52,75,69,67,63,76,72,59,36,
9,7,29,123,170,162,98,31,76,129,149,155,157,159,148,118,83,60,33,20,27,21,21,35,33,37,30,40,36,24,19,24,24,37,54,81,114,77,34,36,43,72,59,47,19,18,23,21,18,16,26,44,65,83,82,90,57,26,72,98,100,98,105,108,111,105,106,108,105,101,101,101,106,111,113,117,123,127,133,137,147,150,159,173,178,186,193,198,201,204,204,219,149,43,52,47,47,52,55,59,68,79,88,107,128,137,124,114,128,195,217,195,127,72,47,45,62,54,44,70,71,66,65,70,78,69,47,27,
14,6,23,123,168,164,115,35,75,128,150,156,157,161,151,110,74,65,32,21,19,17,32,37,27,35,27,40,39,31,22,27,29,27,24,54,96,126,85,71,78,49,17,24,27,20,21,15,15,18,33,55,75,85,88,73,18,45,91,101,100,100,104,106,106,107,109,106,105,104,102,100,104,107,111,115,120,123,129,134,142,147,156,168,175,185,190,196,200,201,204,214,182,58,64,68,60,53,45,38,34,33,34,53,82,117,163,149,151,204,213,170,89,43,29,48,52,48,68,77,62,65,62,74,76,62,35,25,
28,35,39,117,171,174,125,42,76,127,151,157,156,165,154,102,81,54,23,22,25,27,30,30,26,31,31,41,34,33,29,21,23,30,27,20,58,122,122,85,73,71,15,23,19,20,20,16,13,22,43,68,78,85,84,32,21,77,97,101,100,103,104,104,104,108,111,108,107,104,102,101,106,105,107,112,118,122,128,131,136,144,155,165,172,181,189,194,196,202,203,208,207,90,65,78,76,70,59,48,37,22,14,12,41,148,199,153,165,209,205,134,47,27,38,51,42,61,81,69,58,56,67,79,74,52,32,24,
62,60,64,115,168,178,136,57,75,125,152,158,157,166,154,100,86,56,17,25,35,29,21,27,27,28,34,36,41,34,24,21,22,26,42,28,19,64,118,117,79,85,27,21,18,18,15,14,17,37,55,78,87,86,40,18,58,93,98,100,101,106,104,105,105,107,109,111,109,107,105,103,103,105,105,109,113,117,126,128,133,143,151,156,170,179,185,192,198,198,201,204,216,127,56,80,82,77,70,63,52,35,24,9,39,171,197,150,182,206,165,60,22,33,44,41,52,78,74,55,53,56,75,86,68,52,38,31,
63,69,84,126,167,176,147,68,74,126,151,159,160,166,157,97,83,51,22,23,22,23,21,30,28,24,23,37,36,38,36,20,31,37,37,35,39,45,61,90,103,49,20,22,21,18,13,18,30,48,67,87,77,35,15,53,87,93,96,99,103,105,105,105,104,106,110,107,109,107,107,101,102,107,109,108,114,117,121,125,132,140,142,153,164,173,182,190,194,199,201,202,211,167,56,73,83,82,73,67,61,52,39,26,44,150,197,186,181,153,75,21,27,40,36,48,73,76,58,48,50,66,87,80,65,53,36,39,
51,84,95,122,163,170,147,73,76,123,152,157,161,166,156,95,84,42,18,27,28,27,26,30,28,20,31,56,35,50,53,18,30,58,33,49,40,48,79,86,49,49,19,22,20,14,13,25,47,61,63,46,23,27,61,81,90,94,97,101,103,104,104,106,104,107,108,109,113,110,110,108,107,106,104,105,111,114,118,123,131,138,143,147,155,169,176,185,192,196,202,202,208,198,73,64,78,80,76,72,70,59,58,55,61,152,209,189,119,62,30,30,42,39,46,72,80,65,46,47,59,83,85,76,63,42,41,41,
33,71,80,106,157,173,147,78,74,121,151,159,162,166,157,103,65,35,17,28,29,32,27,28,41,21,31,63,39,49,79,36,25,51,23,61,56,36,73,121,56,34,18,20,20,19,19,24,35,28,28,31,50,71,85,89,90,96,96,102,102,102,105,105,104,108,108,112,115,115,113,109,109,106,107,108,108,113,118,123,127,134,139,149,156,163,174,182,189,195,200,203,204,211,106,55,73,77,80,78,77,71,73,74,68,132,177,123,55,45,40,46,45,46,72,87,66,50,38,48,74,89,86,73,49,37,42,35,
25,45,64,93,151,169,149,89,76,118,149,159,162,166,156,113,43,25,22,26,24,35,32,35,46,22,31,57,31,45,95,64,19,62,45,28,72,40,75,102,87,40,21,25,22,18,15,21,29,42,52,68,82,86,90,91,92,93,94,98,100,103,102,102,107,106,107,111,113,114,112,111,113,108,107,110,109,111,116,120,128,132,136,146,156,163,170,178,185,193,196,200,205,213,143,49,67,75,80,86,82,80,89,86,78,89,94,62,52,54,58,50,44,63,81,72,49,38,36,68,88,95,87,68,43,37,34,27,
33,38,48,78,147,181,165,103,79,117,150,159,162,166,157,96,36,34,24,27,22,36,35,33,52,26,28,60,19,40,77,87,18,58,81,16,51,62,49,90,70,42,20,25,18,16,25,44,60,74,76,81,88,90,90,92,95,91,92,99,101,101,100,105,107,107,107,109,112,113,112,114,112,115,113,110,110,114,118,119,123,130,136,142,150,158,166,173,181,187,195,202,200,209,178,54,61,75,81,90,88,92,94,86,83,76,70,64,71,74,60,50,55,72,65,51,46,43,52,83,98,92,79,55,35,31,29,24,
29,30,34,69,167,199,192,130,82,118,151,160,162,167,152,81,32,29,29,21,29,32,31,36,42,37,30,76,18,49,65,93,64,27,77,31,27,75,41,56,75,40,17,18,19,26,43,62,74,81,82,83,88,91,91,91,92,96,95,97,98,100,103,102,102,105,106,107,110,110,114,115,115,116,114,114,115,115,119,122,122,128,136,143,148,156,163,169,178,187,191,198,199,204,199,73,53,74,82,84,94,98,92,86,85,78,75,76,85,79,63,61,73,69,49,42,45,52,75,98,100,84,62,39,31,31,27,33,
27,29,27,69,176,197,195,150,85,117,150,158,158,164,149,95,38,22,27,28,35,34,36,48,37,40,48,74,18,58,63,63,96,16,66,56,29,55,45,36,69,87,49,6,22,40,58,68,74,80,85,84,88,91,89,93,95,95,97,95,98,102,100,99,106,104,104,107,112,113,114,112,115,115,118,117,115,115,121,124,124,126,137,141,144,154,160,170,176,183,191,194,197,203,210,110,48,69,75,82,93,93,94,92,83,83,85,93,91,72,64,69,64,58,57,54,51,71,101,106,90,69,43,28,24,32,43,57,
24,27,24,56,171,194,191,148,86,118,149,160,162,164,150,72,36,20,24,31,31,40,40,47,41,36,87,55,25,57,59,38,76,61,74,58,17,41,47,24,48,56,80,41,39,52,59,70,77,82,86,87,89,95,92,93,93,94,97,93,98,102,101,97,100,103,106,107,112,113,110,111,114,113,119,118,119,119,121,122,130,130,134,141,143,148,155,167,176,181,185,191,196,199,210,147,63,68,67,78,85,93,102,96,90,92,104,104,87,67,59,53,50,60,64,57,61,87,108,105,80,45,26,19,25,44,63,69);
	
	process(blur_matrix_int, blur_matrix)
	begin
		blur_comp14:for i in 0 to matrix_size-1 loop
			blur_comp15:for j in 0 to matrix_size-1 loop
				blur_matrix(i)(j) <= blur_matrix_int((matrix_size*i)+j);
			end loop blur_comp15;
		end loop blur_comp14;

		blur_comp10:for i in 1 to matrix_size-2 loop
			blur_comp11:for j in 1 to matrix_size-2 loop
				blur_sum_matrix(i)(j) <= conv_std_logic_vector((blur_matrix(i-1)(j-1)+blur_matrix(i-1)(j)+blur_matrix(i-1)(j+1)+blur_matrix(i)(j-1)+blur_matrix(i)(j)+blur_matrix(i)(j+1)+blur_matrix(i+1)(j-1)+blur_matrix(i+1)(j)+blur_matrix(i+1)(j+1)),12);
			end loop blur_comp11;
		end loop blur_comp10;
	
		blur_sum_matrix(0)(0) <= conv_std_logic_vector((blur_matrix(0)(0)+blur_matrix(0)(1)+blur_matrix(1)(0)+blur_matrix(1)(1)),12);
		blur_sum_matrix(0)(matrix_size-1) <= conv_std_logic_vector((blur_matrix(0)(matrix_size-2)+blur_matrix(0)(matrix_size-1)+blur_matrix(1)(matrix_size-2)+blur_matrix(1)(matrix_size-1)),12);
		blur_sum_matrix(matrix_size-1)(0) <= conv_std_logic_vector((blur_matrix(matrix_size-2)(0)+blur_matrix(matrix_size-2)(1)+blur_matrix(matrix_size-1)(0)+blur_matrix(matrix_size-1)(1)),12);
		blur_sum_matrix(matrix_size-1)(matrix_size-1) <= conv_std_logic_vector((blur_matrix(matrix_size-2)(matrix_size-2)+blur_matrix(matrix_size-2)(matrix_size-1)+blur_matrix(matrix_size-1)(matrix_size-2)+blur_matrix(matrix_size-1)(matrix_size-1)),12);
		
		blur_comp12:for k in 1 to matrix_size-2 loop
			blur_sum_matrix(0)(k) <= conv_std_logic_vector((blur_matrix(0)(k-1)+blur_matrix(0)(k)+blur_matrix(0)(k+1)+blur_matrix(1)(k-1)+blur_matrix(1)(k)+blur_matrix(1)(k+1)),12);
			blur_sum_matrix(k)(0) <= conv_std_logic_vector((blur_matrix(k-1)(0)+blur_matrix(k-1)(1)+blur_matrix(k)(0)+blur_matrix(k)(1)+blur_matrix(k+1)(0)+blur_matrix(k+1)(1)),12);
			blur_sum_matrix(matrix_size-1)(k) <= conv_std_logic_vector((blur_matrix(matrix_size-2)(k-1)+blur_matrix(matrix_size-2)(k)+blur_matrix(matrix_size-2)(k+1)+blur_matrix(matrix_size-1)(k-1)+blur_matrix(matrix_size-1)(k)+blur_matrix(matrix_size-1)(k+1)),12);
			blur_sum_matrix(k)(matrix_size-1) <= conv_std_logic_vector((blur_matrix(k-1)(matrix_size-2)+blur_matrix(k-1)(matrix_size-1)+blur_matrix(k)(matrix_size-2)+blur_matrix(k)(matrix_size-1)+blur_matrix(k+1)(matrix_size-2)+blur_matrix(k+1)(matrix_size-1)),12);
		end loop blur_comp12;
		
	end process;

	blur_comp0: blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(0)(0),
      							blur_mult_regop2 => "001000000000",
							blur_mult_regres => blur_res_matrix(0)(0));

	blur_comp1: blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(0)(matrix_size-1),
      							blur_mult_regop2 => "001000000000",
							blur_mult_regres => blur_res_matrix(0)(matrix_size-1));
	
	blur_comp2: blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(matrix_size-1)(0),
      							blur_mult_regop2 => "001000000000",
							blur_mult_regres => blur_res_matrix(matrix_size-1)(0));

	blur_comp3: blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(matrix_size-1)(matrix_size-1),
      							blur_mult_regop2 => "001000000000",
							blur_mult_regres => blur_res_matrix(matrix_size-1)(matrix_size-1));
 
	blur_comp4: for m in 1 to matrix_size-2 generate
		blur_comp4_m : blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(0)(m),
      							blur_mult_regop2 => "000101000111",
							blur_mult_regres => blur_res_matrix(0)(m));
	end generate blur_comp4;

	blur_comp5: for m in 1 to matrix_size-2 generate
		blur_comp5_m : blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(m)(0),
      							blur_mult_regop2 => "000101000111",
							blur_mult_regres => blur_res_matrix(m)(0));
	end generate blur_comp5;
	
	blur_comp6: for m in 1 to matrix_size-2 generate
		blur_comp6_m : blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(matrix_size-1)(m),
      							blur_mult_regop2 => "000101000111",
							blur_mult_regres => blur_res_matrix(matrix_size-1)(m));
	end generate blur_comp6;

	blur_comp7: for m in 1 to matrix_size-2 generate
		blur_comp7_m : blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(m)(matrix_size-1),
      							blur_mult_regop2 => "000101000111",
							blur_mult_regres => blur_res_matrix(m)(matrix_size-1));
	end generate blur_comp7;

	blur_comp8: for m in 1 to matrix_size-2 generate
		blur_comp9: for n in 1 to matrix_size-2 generate
			blur_com9_m : blur_mult port map (blur_mult_regxnor_value => blur_xnor_value,
							blur_mult_regop1 => blur_sum_matrix(m)(n),
      							blur_mult_regop2 => "000011100001",
							blur_mult_regres => blur_res_matrix(m)(n));
		end generate blur_comp9;
	end generate blur_comp8;
	

	process
	variable l: line;
	file outfile: text open write_mode is "C:\Modeltech_pe_edu_10.4a\examples\output.txt";
	begin
		wait for 9999 ns;
		blur_comp16: for p in 0 to matrix_size-1 loop
			blur_comp17: for q in 0 to matrix_size-1 loop
				write(l, blur_res_matrix(p)(q));
				writeline(outfile, l);
			end loop blur_comp17;
		end loop blur_comp16;
	end process;


end blur_arch;
