library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.math_real.all;
use IEEE.STD_LOGIC_TEXTIO.ALL;
use STD.TEXTIO.ALL;

library work;
use work.blur_pkg.all;

entity tb_blur is
end tb_blur;


architecture tb_blur_behav of tb_blur is

component blur is
port
   (
	blur_clk : in std_logic;
	blur_xnor_value : in std_logic_vector (12 downto 0);
	blur_matrix_int : in blur_matrix_int_type;
	blur_res_matrix : out blur_res_matrix_type
   );
end component;
  
signal t_blur_clk : std_logic := '0';
signal t_blur_xnor_value : std_logic_vector (12 downto 0);
signal t_blur_matrix_int : blur_matrix_int_type;
signal t_blur_res_matrix : blur_res_matrix_type;


begin

	U1 : blur port map (t_blur_clk, t_blur_xnor_value, t_blur_matrix_int, t_blur_res_matrix);
	t_blur_clk <= not (t_blur_clk) after 5 ns;
	--clk_process :process
   	--begin
        	--t_blur_clk <= '0';
        	--wait for 5 ns;
        	--t_blur_clk <= '1';
        	--wait for 5 ns;
   	--end process;

	test_process : process
	begin
		wait until t_blur_clk = '1' and t_blur_clk'event;
		t_blur_xnor_value <= "0000000000000";
		t_blur_matrix_int <= (137,135,133,136,138,133,135,132,137,137,133,136,137,135,134,132,138,133,134,135,136,131,130,130,133,133,132,130,134,133,128,125,129,132,131,130,134,131,132,128,131,134,130,122,132,130,130,130,131,130,130,130,132,132,127,130,131,132,130,130,131,131,131,128);
		wait for 10 ns;
		t_blur_matrix_int <= (132,139,129,130,132,127,129,129,132,138,130,131,132,127,129,129,131,134,127,127,131,127,128,130,129,128,129,124,128,127,123,131,127,132,129,126,130,126,126,130,131,127,132,128,124,128,129,126,130,131,133,128,127,128,127,129,129,129,128,128,128,127,127,131);
		wait for 10 ns;
		t_blur_matrix_int <= (131,130,139,138,142,146,151,151,130,131,138,138,142,147,151,151,130,128,136,138,143,145,150,150,131,128,132,140,144,146,149,149,126,132,137,143,146,146,147,149,128,131,138,143,145,146,150,147,131,139,140,145,147,147,145,146,136,142,144,146,146,146,146,144);
		wait for 10 ns;
		t_blur_matrix_int <= (148,149,142,134,119,118,90,80,150,147,143,134,119,118,91,79,148,149,143,133,119,110,88,78,150,146,141,130,120,102,90,76,149,145,140,127,116,106,87,78,148,144,142,124,110,102,91,74,145,141,140,125,112,103,85,73,142,141,130,127,113,98,87,78);
		wait for 10 ns;
		t_blur_matrix_int <= (64,62,60,70,70,73,73,74,65,61,61,68,72,72,73,74,65,60,61,65,69,68,73,75,60,55,57,60,62,65,74,76,61,57,55,57,64,67,67,69,59,56,55,60,64,65,64,71,63,55,57,61,59,65,67,73,62,60,59,60,62,70,67,69);
		wait for 10 ns;
		t_blur_matrix_int <= (78,74,76,79,76,75,78,76,78,75,76,78,76,75,78,76,76,73,73,76,72,73,77,73,68,71,69,72,70,72,73,72,72,70,67,75,72,74,73,71,65,72,69,72,72,72,67,71,70,74,74,77,77,71,66,73,72,74,76,73,74,70,68,72);
		wait for 10 ns;
		t_blur_matrix_int <= (78,78,74,74,79,83,83,88,78,78,74,74,80,82,83,88,76,76,74,75,78,80,83,87,70,73,72,74,76,79,86,85,71,72,74,75,79,79,80,84,73,68,72,75,78,79,80,86,68,69,69,74,82,79,82,86,75,66,68,74,78,77,80,84);
		wait for 10 ns;
		t_blur_matrix_int <= (84,90,93,91,95,94,91,102,83,90,93,92,96,93,91,102,86,89,92,91,93,94,90,97,86,92,94,93,93,89,91,94,84,89,88,92,93,93,92,98,87,90,92,93,90,93,90,98,86,85,89,88,93,92,93,91,84,86,91,93,94,93,93,98);
		wait for 10 ns;
		t_blur_matrix_int <= (97,101,97,97,107,102,100,97,98,101,97,97,107,102,101,96,99,100,99,97,105,99,100,100,98,95,101,96,97,100,97,96,91,95,94,99,99,97,97,99,93,98,95,96,96,96,94,101,93,91,94,97,96,97,99,101,94,94,97,94,94,96,99,99);
		wait for 10 ns;
		t_blur_matrix_int <= (97,96,103,99,99,97,105,104,97,95,103,98,100,98,103,104,97,98,101,100,97,98,104,103,98,102,99,99,99,97,98,97,99,96,99,97,100,98,99,102,100,99,101,97,100,97,95,102,99,100,97,97,97,97,99,100,97,99,97,97,98,95,98,99);
		wait for 10 ns;
		t_blur_matrix_int <= (98,101,102,103,101,101,101,101,98,101,102,103,102,101,101,101,100,104,103,104,100,102,102,101,99,100,102,102,101,97,101,101,98,100,101,102,101,104,103,99,96,100,102,103,97,98,99,100,95,98,103,97,98,99,103,103,99,99,98,96,97,102,99,99);
		wait for 10 ns;
		t_blur_matrix_int <= (103,103,101,100,101,106,101,101,103,103,102,100,103,104,101,101,102,106,100,98,100,102,100,100,100,96,102,98,97,99,97,100,98,103,103,100,98,106,102,99,100,100,99,94,97,102,97,100,98,97,98,103,100,100,99,98,98,97,99,99,100,101,99,96);
		wait for 10 ns;
		t_blur_matrix_int <= (105,102,106,104,105,103,104,104,105,103,104,106,105,103,104,103,104,101,103,101,104,103,102,103,101,102,100,101,101,100,98,99,102,99,96,100,98,100,98,95,100,97,99,102,97,99,99,98,95,99,95,100,95,98,98,101,95,101,100,102,99,101,96,98);
		wait for 10 ns;
		t_blur_matrix_int <= (107,104,102,101,100,101,101,99,107,104,102,101,100,101,101,99,103,106,101,98,97,100,100,98,106,100,108,97,105,97,100,96,96,99,98,103,97,96,93,96,97,100,99,98,98,100,96,97,99,100,99,99,97,95,98,94,99,100,99,98,99,98,98,100);
		wait for 10 ns;
		t_blur_matrix_int <= (99,106,105,100,100,100,97,101,99,106,105,100,100,100,97,101,99,102,106,98,98,100,96,102,98,106,105,97,102,93,99,100,102,102,104,100,92,95,98,100,96,96,100,98,99,98,98,97,97,99,99,99,95,95,100,98,99,100,99,99,94,99,100,98);
		wait for 10 ns;
		t_blur_matrix_int <= (104,102,103,106,100,102,97,105,104,102,103,105,101,102,96,105,101,102,102,103,100,100,97,103,103,101,101,98,101,96,101,99,99,97,97,99,97,97,98,99,100,98,103,99,99,96,96,97,103,103,103,100,101,99,100,98,99,103,100,103,101,96,102,98);
		wait for 10 ns;
		t_blur_matrix_int <= (111,103,99,97,101,98,103,98,111,103,98,98,101,99,101,98,106,103,99,98,98,99,98,99,102,102,99,97,95,96,95,101,99,101,100,96,97,97,94,99,96,97,100,99,98,97,96,96,98,100,97,98,103,99,95,99,96,100,100,98,96,98,100,98);
		wait for 10 ns;
		t_blur_matrix_int <= (98,101,96,106,98,99,98,98,98,101,96,105,98,99,98,99,97,99,97,105,93,97,99,100,93,97,98,95,95,97,98,97,92,97,96,95,92,94,92,93,96,96,97,97,95,97,96,97,94,98,97,97,94,98,95,98,97,95,96,94,96,96,95,98);
		wait for 10 ns;
		t_blur_matrix_int <= (99,97,97,97,99,94,99,98,99,97,97,97,98,94,98,98,96,97,97,97,98,95,95,97,98,97,96,95,96,95,94,94,98,97,93,96,98,91,93,94,94,96,100,95,96,97,97,95,94,93,95,97,94,96,101,94,95,96,98,96,96,100,96,94);
		wait for 10 ns;
		t_blur_matrix_int <= (92,91,90,90,87,84,80,72,92,91,89,89,88,84,79,72,92,90,91,90,85,83,79,74,91,89,92,87,84,83,75,75,94,92,88,87,83,79,81,76,93,93,85,90,83,85,77,77,92,91,92,89,85,79,80,82,94,93,91,88,88,80,83,86);
		wait for 10 ns;
		t_blur_matrix_int <= (76,85,96,108,113,121,128,130,76,85,96,108,113,121,127,131,74,84,95,106,111,121,126,129,69,83,91,99,108,119,123,129,71,74,82,93,101,112,120,123,75,72,76,87,100,107,114,121,80,72,72,82,95,106,113,118,78,74,73,78,86,100,111,118);
		wait for 10 ns;
		t_blur_matrix_int <= (136,138,141,131,121,125,126,127,136,138,140,130,120,125,128,127,134,138,138,131,125,127,126,126,133,135,135,131,128,126,125,127,129,131,139,132,130,130,127,126,125,133,135,133,131,128,131,127,125,127,134,136,135,133,130,133,122,126,132,137,136,137,135,136);
		wait for 10 ns;
		t_blur_matrix_int <= (128,127,129,128,134,130,128,128,129,127,131,127,134,130,128,128,124,127,130,127,130,131,128,127,125,127,127,126,128,130,127,127,131,131,130,128,132,128,129,130,129,132,133,132,133,129,131,131,129,134,134,136,136,137,134,132,133,135,137,138,138,139,136,132);
		wait for 10 ns;
		t_blur_matrix_int <= (126,126,127,127,125,130,130,127,126,128,126,127,125,130,128,127,127,125,126,128,127,127,133,128,129,126,127,127,130,127,128,125,131,129,128,126,127,129,125,129,132,129,128,129,128,132,129,127,131,131,129,130,132,131,130,128,132,130,128,129,129,130,126,130);
		wait for 10 ns;
		t_blur_matrix_int <= (130,132,134,129,133,136,132,128,131,132,134,129,134,137,131,129,131,129,133,130,132,133,133,128,127,130,130,130,131,133,128,130,129,132,129,128,128,128,128,129,127,129,124,128,128,131,127,127,129,126,130,127,125,130,128,128,129,130,125,123,125,126,128,127);
		wait for 10 ns;
		t_blur_matrix_int <= (133,147,185,199,206,208,212,212,132,148,184,200,205,207,212,211,129,144,182,198,204,208,211,211,126,130,161,189,201,207,210,212,129,125,136,174,194,203,208,211,130,123,126,151,184,198,206,209,130,124,125,132,168,191,201,207,126,129,126,121,147,182,196,205);
		wait for 10 ns;
		t_blur_matrix_int <= (212,201,168,113,77,72,79,79,212,200,170,113,76,73,79,79,213,203,176,122,77,71,75,82,213,210,195,157,100,71,73,79,210,212,206,183,132,83,77,77,210,213,211,198,163,108,73,73,211,213,213,209,187,142,87,75,210,213,213,213,201,175,123,76);
		wait for 10 ns;
		t_blur_matrix_int <= (88,89,90,93,98,88,93,89,87,90,89,94,98,87,94,89,89,88,89,92,94,90,92,90,85,85,90,83,91,89,90,95,82,82,87,90,91,90,89,93,76,81,83,85,91,90,88,93,77,84,84,83,87,89,88,92,77,77,77,79,89,83,86,91);
		wait for 10 ns;
		t_blur_matrix_int <= (93,99,91,92,90,91,90,90,93,99,91,93,90,91,90,89,94,97,91,90,90,89,90,92,90,95,92,94,95,92,94,96,91,93,91,93,87,90,92,94,89,92,90,91,90,90,88,92,92,90,90,91,89,87,93,91,88,89,96,90,87,92,89,91);
		wait for 10 ns;
		t_blur_matrix_int <= (94,93,95,95,96,93,94,86,94,92,96,95,95,94,94,86,94,94,93,94,96,95,93,87,95,95,96,93,92,92,91,94,95,91,95,90,95,92,94,93,90,93,92,94,93,91,93,91,94,92,93,88,94,91,92,90,91,89,91,93,93,95,94,93);
		wait for 10 ns;
		t_blur_matrix_int <= (97,95,98,96,91,99,96,91,96,96,99,96,91,98,98,90,96,93,98,95,94,99,95,91,89,94,96,91,92,97,97,94,92,96,96,96,95,96,97,99,93,93,93,94,92,95,100,102,97,95,92,96,93,93,105,103,93,95,95,98,100,102,106,90);
		wait for 10 ns;
		t_blur_matrix_int <= (85,86,85,92,123,145,147,114,86,85,86,92,123,144,148,114,85,87,89,93,116,133,125,87,91,91,96,99,85,69,44,30,97,94,95,78,47,28,22,20,103,95,72,43,24,21,21,24,92,79,42,37,19,18,22,24,69,37,22,29,24,22,26,26);
		wait for 10 ns;
		t_blur_matrix_int <= (129,129,130,127,130,129,130,129,129,131,132,129,131,129,132,134,130,130,128,129,131,130,133,132,131,129,126,130,132,130,131,132,129,128,127,130,132,132,132,132,128,130,129,129,131,133,133,130,130,133,132,132,131,131,133,132,131,133,132,132,133,132,136,135);
		wait for 10 ns;
		t_blur_matrix_int <= (127,129,130,129,124,126,128,138,134,134,128,130,129,129,132,137,133,131,127,128,127,130,133,140,134,131,131,133,127,128,131,136,136,129,131,132,129,134,136,142,133,134,129,131,132,136,141,142,132,134,132,133,135,141,144,147,135,134,135,139,140,143,143,147);
		wait for 10 ns;
		t_blur_matrix_int <= (138,144,145,144,145,141,143,141,141,143,144,144,145,142,142,138,141,144,139,145,142,140,141,137,145,147,144,139,143,141,140,137,143,143,146,143,139,138,138,130,143,145,142,144,136,135,135,135,148,145,144,139,134,135,132,134,146,144,142,137,134,133,129,135);
		wait for 10 ns;
		t_blur_matrix_int <= (142,137,131,124,111,102,87,72,142,135,130,121,113,107,93,80,137,137,130,125,113,102,95,85,133,137,130,123,118,104,97,79,135,135,131,125,116,103,88,76,135,134,136,125,116,102,84,69,138,137,134,127,115,103,87,73,135,137,137,128,114,101,89,75);
		wait for 10 ns;
		t_blur_matrix_int <= (59,55,54,59,57,70,70,63,64,56,56,62,62,67,66,66,66,61,56,60,62,65,69,69,63,56,59,62,66,65,67,69,63,54,54,62,60,60,66,74,55,57,47,54,61,65,68,70,60,52,52,59,65,63,68,71,60,57,51,59,64,65,66,69);
		wait for 10 ns;
		t_blur_matrix_int <= (74,72,72,77,71,70,71,73,70,70,77,71,71,72,72,70,78,73,70,75,70,73,67,67,81,68,69,68,68,72,70,71,73,72,72,66,75,74,69,69,68,71,73,76,72,73,68,70,68,72,72,71,75,70,75,70,75,76,77,68,76,70,69,70);
		wait for 10 ns;
		t_blur_matrix_int <= (68,68,67,69,77,78,81,81,68,73,69,75,77,82,84,82,76,68,68,70,79,78,81,81,69,74,72,71,76,80,77,84,70,68,70,76,75,81,75,81,69,68,71,73,77,72,81,82,73,68,72,75,74,75,82,83,73,68,72,73,74,75,78,83);
		wait for 10 ns;
		t_blur_matrix_int <= (83,87,89,91,92,91,93,95,90,87,88,87,93,91,89,95,85,86,87,91,92,89,90,93,83,89,87,87,90,91,91,91,87,90,88,87,91,87,96,94,87,89,85,90,90,93,88,97,83,87,89,89,89,92,92,96,84,87,91,90,91,92,92,90);
		wait for 10 ns;
		t_blur_matrix_int <= (96,94,95,100,95,96,99,98,96,93,95,97,94,97,100,99,92,95,96,96,96,96,99,96,94,95,95,99,98,95,99,94,94,96,91,92,98,98,96,98,95,97,94,93,93,94,96,97,95,95,92,93,95,94,96,95,95,92,95,94,96,95,95,93);
		wait for 10 ns;
		t_blur_matrix_int <= (97,98,98,98,102,97,95,97,99,98,102,99,100,98,97,100,95,101,94,98,99,99,98,100,99,98,100,96,95,97,96,98,94,96,97,97,94,95,97,96,94,95,95,95,95,98,97,99,92,97,95,96,97,100,92,98,94,92,96,95,96,97,97,95);
		wait for 10 ns;
		t_blur_matrix_int <= (99,102,101,100,98,103,102,100,97,98,99,95,97,100,100,99,98,96,99,100,97,97,98,99,96,99,100,97,98,98,99,97,95,96,98,96,94,98,101,100,97,100,96,94,91,98,94,96,97,98,97,99,97,95,95,100,95,101,94,99,98,96,96,98);
		wait for 10 ns;
		t_blur_matrix_int <= (106,101,101,97,100,101,101,99,99,102,98,97,98,99,98,97,100,95,97,99,95,98,98,99,98,95,99,96,97,94,99,96,95,97,94,96,94,96,98,102,96,97,94,93,96,99,98,99,93,97,91,93,94,93,95,101,94,97,96,95,94,95,98,100);
		wait for 10 ns;
		t_blur_matrix_int <= (97,96,101,101,100,96,101,102,98,93,98,107,99,99,100,99,98,96,101,98,97,95,94,101,98,100,93,97,99,91,95,98,103,100,96,96,94,94,93,93,103,102,101,96,93,88,89,91,102,104,102,97,91,90,91,91,100,96,98,99,95,95,88,90);
		wait for 10 ns;
		t_blur_matrix_int <= (101,103,101,98,102,100,96,95,97,97,100,99,103,98,99,98,101,97,97,97,98,98,106,98,93,94,94,97,96,96,92,98,90,93,93,90,94,93,92,94,90,90,90,92,91,97,94,95,89,86,87,90,86,92,98,94,84,88,90,88,91,90,91,95);
		wait for 10 ns;
		t_blur_matrix_int <= (95,102,100,99,98,95,98,100,95,103,103,101,95,95,97,99,101,99,99,98,94,95,98,97,98,97,96,99,94,95,95,97,92,94,93,94,94,95,92,93,95,91,92,94,95,93,93,98,91,92,91,91,89,93,94,93,93,93,92,91,93,90,92,93);
		wait for 10 ns;
		t_blur_matrix_int <= (102,104,103,106,101,99,100,97,102,102,104,106,102,99,101,100,99,101,103,106,111,101,100,96,102,98,100,101,102,98,98,97,97,97,97,101,99,99,98,99,90,96,93,97,102,98,99,98,95,98,98,94,97,96,98,98,91,99,99,96,95,99,98,100);
		wait for 10 ns;
		t_blur_matrix_int <= (101,98,99,97,100,98,94,96,101,99,97,103,101,96,96,92,101,97,98,98,102,96,97,94,96,97,99,97,98,101,96,96,98,99,98,100,95,96,93,92,100,100,97,103,94,94,94,95,98,99,104,98,97,92,95,93,101,96,100,92,97,93,97,92);
		wait for 10 ns;
		t_blur_matrix_int <= (97,96,96,96,93,91,95,95,97,99,99,98,96,95,93,96,97,95,96,96,96,91,90,95,96,99,90,92,93,92,94,95,94,96,97,92,94,91,91,93,93,95,92,93,97,93,93,96,95,95,97,96,94,92,96,91,92,98,94,95,98,92,90,94);
		wait for 10 ns;
		t_blur_matrix_int <= (98,98,98,96,98,95,97,97,96,96,99,98,97,91,96,97,95,94,96,96,94,95,95,94,93,96,92,94,89,92,97,96,95,96,93,92,91,91,96,95,96,94,95,91,93,98,94,93,92,92,93,91,89,97,94,95,95,90,93,92,93,98,94,96);
		wait for 10 ns;
		t_blur_matrix_int <= (95,96,89,89,84,81,84,89,94,98,93,90,86,83,83,80,94,91,94,90,102,86,81,83,92,92,90,91,88,89,81,81,92,91,94,90,95,85,82,77,92,94,89,91,94,94,81,77,92,90,94,85,86,87,88,79,96,98,87,84,86,85,86,83);
		wait for 10 ns;
		t_blur_matrix_int <= (77,79,74,71,82,94,111,117,78,77,71,69,81,90,101,111,77,74,77,70,78,87,100,111,79,83,74,74,78,80,96,106,77,76,75,76,84,89,97,107,78,77,72,74,80,88,91,102,81,77,76,76,80,87,96,101,76,78,78,74,79,91,99,104);
		wait for 10 ns;
		t_blur_matrix_int <= (118,125,131,132,136,142,137,135,120,126,130,132,136,138,137,138,121,122,128,131,137,139,139,141,119,122,128,132,136,137,138,138,116,123,126,133,136,137,139,137,110,118,127,134,133,135,137,135,113,117,126,130,131,133,136,139,107,118,123,127,132,129,133,139);
		wait for 10 ns;
		t_blur_matrix_int <= (134,134,137,139,135,139,137,133,137,134,137,138,141,136,140,139,137,134,136,137,136,141,135,136,134,138,135,136,135,141,135,136,140,141,134,134,136,136,135,136,137,135,136,134,133,135,133,134,137,135,137,134,135,135,136,130,134,135,132,130,133,132,136,133);
		wait for 10 ns;
		t_blur_matrix_int <= (132,133,137,134,131,128,127,126,133,132,133,134,134,131,130,127,136,131,131,130,131,131,127,130,138,137,131,128,130,130,127,128,134,137,132,127,129,132,129,129,135,135,135,131,130,132,130,131,136,133,132,133,132,129,131,129,133,131,132,131,131,128,129,129);
		wait for 10 ns;
		t_blur_matrix_int <= (124,128,132,124,126,123,128,125,128,129,129,125,127,126,125,127,129,131,125,127,125,127,128,129,126,128,125,127,124,126,125,125,129,128,127,127,126,127,124,125,130,128,128,127,127,128,127,125,131,127,131,130,129,132,127,125,131,128,125,131,132,131,129,130);
		wait for 10 ns;
		t_blur_matrix_int <= (126,125,124,122,127,165,190,202,127,127,124,123,120,136,176,196,126,124,124,124,124,120,155,187,124,123,124,126,117,118,133,171,127,125,124,123,121,120,120,150,128,124,126,126,119,121,118,127,127,125,127,123,120,120,120,118,126,127,122,127,121,118,119,116);
		wait for 10 ns;
		t_blur_matrix_int <= (208,211,214,213,210,194,157,98,206,211,213,213,212,204,180,132,201,207,210,213,215,211,198,166,195,204,209,212,214,215,209,188,185,199,208,212,213,216,215,202,171,195,203,210,214,216,217,212,143,183,200,207,211,213,216,216,123,166,191,203,209,213,217,217);
		wait for 10 ns;
		t_blur_matrix_int <= (73,76,78,80,88,83,86,89,78,73,77,79,83,86,83,87,105,75,81,78,85,79,88,87,139,85,74,81,80,82,86,89,175,119,74,73,80,83,87,93,194,156,91,75,78,82,86,82,208,184,129,73,77,79,83,85,215,202,166,101,73,79,79,85);
		wait for 10 ns;
		t_blur_matrix_int <= (89,91,92,89,91,95,91,94,89,92,94,91,95,97,92,93,88,89,92,96,90,90,92,96,87,85,86,90,95,91,92,88,89,92,90,93,93,90,93,89,97,93,96,89,94,94,90,92,86,90,91,94,92,91,92,89,85,88,85,94,93,89,90,91);
		wait for 10 ns;
		t_blur_matrix_int <= (93,94,96,95,92,98,96,96,94,96,94,95,94,97,96,94,90,94,95,105,96,97,98,101,92,89,97,97,101,100,100,100,90,89,94,98,92,99,101,100,86,97,94,91,96,98,100,103,91,91,92,98,93,101,101,106,94,95,91,95,98,103,102,89);
		wait for 10 ns;
		t_blur_matrix_int <= (98,98,97,99,103,103,92,64,98,100,102,102,105,88,62,35,100,104,105,107,92,64,35,22,102,105,107,92,62,30,30,21,105,105,93,59,35,53,25,18,105,94,61,28,19,26,24,15,90,56,26,14,14,22,20,22,60,22,13,20,21,19,23,18);
		wait for 10 ns;
		t_blur_matrix_int <= (32,21,19,18,24,24,14,24,16,23,25,18,27,21,19,22,20,30,28,23,21,24,23,24,27,26,32,23,21,23,24,28,21,19,18,20,20,24,28,29,14,18,19,22,16,27,28,19,18,21,23,22,23,26,23,38,25,20,22,23,23,20,29,30);
		wait for 10 ns;
		t_blur_matrix_int <= (129,131,132,128,133,133,134,134,135,133,133,131,133,137,137,135,133,133,132,135,138,141,135,137,137,135,136,134,134,135,134,137,138,138,138,135,134,139,137,138,133,135,137,135,134,136,135,143,137,132,138,135,136,134,139,146,139,137,137,134,133,139,139,145);
		wait for 10 ns;
		t_blur_matrix_int <= (135,137,134,139,144,147,148,147,135,138,140,141,146,144,144,144,139,140,144,146,145,144,144,145,140,143,145,144,142,142,141,137,141,145,146,142,142,135,136,140,144,147,143,136,136,134,132,134,150,146,138,132,128,130,127,130,144,136,134,128,124,125,120,122);
		wait for 10 ns;
		t_blur_matrix_int <= (146,144,144,137,136,134,132,134,143,142,145,135,134,134,133,133,144,141,138,133,130,132,134,133,139,140,136,135,131,133,136,135,139,136,136,133,134,133,135,135,132,130,135,135,134,132,134,134,128,130,135,139,136,135,133,133,124,127,136,138,140,137,132,139);
		wait for 10 ns;
		t_blur_matrix_int <= (136,136,134,126,118,104,91,72,135,139,134,125,114,101,84,72,134,134,133,124,112,100,92,72,135,136,132,125,112,104,87,70,136,135,130,126,111,98,86,65,134,137,134,122,112,103,89,69,138,137,133,123,117,98,87,68,137,136,131,127,116,105,91,71);
		wait for 10 ns;
		t_blur_matrix_int <= (60,57,58,63,62,65,64,68,61,54,59,59,64,64,65,72,60,52,53,57,65,62,65,69,54,47,49,56,62,66,67,68,58,46,50,60,56,66,71,73,55,49,51,57,59,67,68,69,61,47,51,61,61,65,67,68,58,51,50,59,60,61,67,69);
		wait for 10 ns;
		t_blur_matrix_int <= (70,72,76,75,78,70,66,67,71,71,72,74,70,70,72,69,70,68,68,69,71,72,68,68,71,74,67,71,70,67,71,71,70,65,66,67,69,69,69,69,67,72,72,71,71,75,64,73,69,68,71,69,65,73,71,69,70,71,74,76,71,69,70,70);
		wait for 10 ns;
		t_blur_matrix_int <= (68,68,71,70,74,77,79,80,67,66,67,69,76,80,78,82,66,73,73,69,77,77,81,80,71,70,66,69,76,78,82,82,67,69,71,69,70,77,79,82,67,67,72,69,73,75,77,81,70,70,69,71,75,74,79,84,69,69,71,70,79,77,82,81);
		wait for 10 ns;
		t_blur_matrix_int <= (84,83,89,91,92,86,91,92,83,84,87,86,90,89,93,91,87,82,88,86,85,87,94,90,83,83,89,85,86,87,86,94,84,88,86,89,88,91,91,87,84,88,89,85,84,89,92,91,82,84,87,86,88,92,93,90,84,87,86,90,85,90,89,89);
		wait for 10 ns;
		t_blur_matrix_int <= (94,94,98,90,95,94,97,94,91,92,95,94,94,93,94,96,86,94,96,94,93,91,99,94,92,91,92,95,92,93,95,93,93,87,88,93,92,92,93,94,92,88,88,89,90,92,96,88,92,94,92,91,92,94,89,91,91,89,91,93,91,92,93,91);
		wait for 10 ns;
		t_blur_matrix_int <= (93,93,93,96,96,95,96,96,94,96,90,93,88,94,95,99,92,92,87,95,87,93,92,96,93,90,87,92,95,95,93,95,91,90,88,90,88,91,92,91,91,91,87,94,94,96,93,94,89,92,94,93,93,94,98,91,91,93,94,97,92,90,95,94);
		wait for 10 ns;
		t_blur_matrix_int <= (95,95,96,97,99,97,98,95,97,94,94,91,94,99,94,96,93,91,96,92,94,91,94,95,96,93,96,93,90,96,96,95,94,94,94,92,91,97,95,93,92,91,92,92,90,95,90,95,94,92,90,91,95,98,95,94,95,93,90,92,92,107,93,96);
		wait for 10 ns;
		t_blur_matrix_int <= (95,97,101,96,93,94,96,95,95,94,95,96,93,96,93,97,95,97,103,97,95,95,95,91,93,96,96,96,96,94,92,94,96,93,95,92,96,95,91,93,95,92,94,95,95,91,95,94,94,97,92,97,90,94,89,91,98,101,92,92,93,88,95,90);
		wait for 10 ns;
		t_blur_matrix_int <= (99,98,98,92,92,97,91,87,98,100,97,94,94,91,90,86,95,95,92,93,88,92,91,90,98,91,93,92,90,90,90,89,94,94,93,92,92,93,93,91,95,92,92,94,89,92,99,93,98,99,90,94,88,89,90,94,94,104,95,90,91,91,98,94);
		wait for 10 ns;
		t_blur_matrix_int <= (89,90,87,86,90,86,91,93,88,90,88,87,87,88,90,92,92,91,88,89,92,89,95,93,92,89,83,92,88,86,87,90,92,90,88,92,88,89,83,85,89,91,90,91,87,89,88,86,91,89,88,89,88,100,102,136,120,113,116,115,120,132,158,148);
		wait for 10 ns;
		t_blur_matrix_int <= (93,90,93,92,92,90,91,92,94,97,89,91,87,89,90,93,93,92,87,88,92,88,85,93,90,85,86,83,86,83,90,89,87,86,87,88,87,86,87,86,84,87,85,87,83,86,84,88,117,134,120,118,104,107,89,88,159,156,161,154,168,164,162,158);
		wait for 10 ns;
		t_blur_matrix_int <= (90,94,98,94,98,96,93,96,90,95,96,97,95,101,97,97,90,92,96,96,97,96,101,97,91,92,90,96,93,94,98,97,87,87,95,95,92,98,101,96,85,86,91,90,93,92,94,96,86,87,88,90,88,87,95,91,128,116,89,87,81,84,86,87);
		wait for 10 ns;
		t_blur_matrix_int <= (103,97,99,95,95,94,94,94,101,102,102,97,94,98,94,96,100,98,102,97,97,93,94,94,101,97,97,94,93,93,94,93,98,96,95,94,93,95,89,94,97,98,95,91,93,94,94,95,90,92,88,94,94,94,94,94,87,92,89,90,89,92,88,95);
		wait for 10 ns;
		t_blur_matrix_int <= (97,97,94,94,96,94,89,95,97,96,92,93,93,93,93,93,95,97,95,93,93,93,89,89,94,96,96,89,93,96,91,93,93,94,96,93,92,88,93,94,88,96,97,101,90,92,96,94,93,94,97,97,95,92,94,92,92,97,98,96,98,95,94,89);
		wait for 10 ns;
		t_blur_matrix_int <= (95,91,92,90,94,92,94,95,93,91,92,92,94,93,93,95,90,94,94,90,92,92,92,93,93,90,91,92,95,91,91,93,95,93,93,93,92,92,94,92,92,94,91,92,88,94,93,94,92,96,98,91,93,93,93,93,91,93,91,90,88,95,91,91);
		wait for 10 ns;
		t_blur_matrix_int <= (93,94,91,87,87,84,82,81,95,93,91,87,87,82,85,79,95,86,86,89,87,81,87,83,93,88,91,86,83,86,87,87,92,91,89,84,85,82,83,82,89,89,89,87,81,87,82,83,92,89,94,88,83,82,82,82,90,90,87,86,83,82,80,83);
		wait for 10 ns;
		t_blur_matrix_int <= (76,76,71,73,76,88,94,100,81,80,74,76,81,86,89,97,84,80,73,73,78,85,91,98,85,77,73,72,75,83,91,100,81,80,79,76,78,84,90,97,80,82,79,74,77,82,87,91,86,79,74,73,76,79,83,93,82,76,75,72,77,84,85,95);
		wait for 10 ns;
		t_blur_matrix_int <= (106,112,119,124,128,131,134,134,104,112,119,124,124,129,130,133,105,110,115,122,126,128,130,128,103,111,119,122,120,127,127,128,102,111,114,119,119,124,126,127,105,107,112,117,120,121,122,126,104,108,111,118,117,119,121,125,102,107,113,115,116,115,117,120);
		wait for 10 ns;
		t_blur_matrix_int <= (135,137,132,135,133,133,135,136,132,135,133,130,133,132,134,133,131,132,130,134,129,133,133,134,131,131,133,133,130,134,129,131,127,130,129,133,132,129,132,130,128,125,132,130,132,126,130,128,124,124,128,129,130,132,128,127,123,122,128,128,127,131,128,130);
		wait for 10 ns;
		t_blur_matrix_int <= (132,135,133,132,132,131,130,131,132,131,130,131,134,133,129,130,133,129,132,128,134,131,127,132,130,131,128,129,132,129,125,126,129,128,130,129,130,127,126,125,127,130,128,129,127,126,127,129,127,128,129,126,129,128,127,130,125,125,126,125,127,127,129,127);
		wait for 10 ns;
		t_blur_matrix_int <= (131,128,131,128,134,130,130,131,131,132,128,127,129,128,130,130,131,130,131,128,131,131,128,127,129,133,131,132,128,130,127,126,127,130,133,130,129,128,128,125,126,127,125,129,127,126,126,124,128,125,127,128,127,125,122,122,127,128,123,125,124,124,121,117);
		wait for 10 ns;
		t_blur_matrix_int <= (128,128,126,126,126,123,118,114,130,125,127,125,126,120,121,115,131,125,124,123,123,120,124,118,126,127,121,121,122,122,119,117,125,125,122,123,123,117,117,115,122,119,121,117,115,119,114,116,121,119,117,113,121,112,113,116,120,118,119,117,117,114,115,117);
		wait for 10 ns;
		t_blur_matrix_int <= (111,130,172,196,204,211,215,218,116,118,159,191,202,211,215,218,116,114,129,172,198,207,214,216,113,112,113,149,188,202,212,217,116,111,110,126,173,199,208,215,112,113,110,115,147,187,204,213,113,114,112,114,124,168,197,206,112,118,115,112,112,141,182,199);
		wait for 10 ns;
		t_blur_matrix_int <= (219,214,198,154,91,77,77,80,220,218,205,179,118,75,72,78,217,219,213,197,158,94,68,69,217,219,219,210,190,131,74,68,218,220,221,216,201,169,102,69,216,218,218,220,210,189,138,77,213,218,218,219,218,203,172,104,211,215,218,219,219,212,195,149);
		wait for 10 ns;
		t_blur_matrix_int <= (85,87,85,87,89,95,94,93,80,81,87,85,92,93,89,91,79,82,83,83,89,94,93,97,79,78,80,82,85,87,88,95,75,79,76,80,82,83,91,92,71,76,76,79,80,82,89,92,70,74,74,80,85,81,94,98,82,87,79,82,85,89,95,85);
		wait for 10 ns;
		t_blur_matrix_int <= (97,92,95,99,103,102,91,66,92,101,98,100,103,93,61,27,95,101,101,101,86,58,28,15,97,100,104,88,62,27,17,21,100,98,91,63,29,20,17,20,104,89,61,33,19,17,14,18,88,63,30,21,19,18,19,20,55,31,20,18,21,24,18,21);
		wait for 10 ns;
		t_blur_matrix_int <= (35,13,21,13,30,26,25,17,17,14,15,18,22,33,25,28,17,15,20,24,25,26,28,28,19,19,15,27,34,39,33,36,16,20,20,25,25,27,28,25,21,21,28,30,34,37,30,25,22,24,26,30,31,34,30,29,22,25,28,31,33,35,31,28);
		wait for 10 ns;
		t_blur_matrix_int <= (28,25,26,22,23,23,29,32,27,18,26,22,23,29,27,21,24,25,26,22,21,29,21,19,35,26,26,26,22,19,19,26,24,26,20,19,22,18,19,20,28,26,24,23,18,18,20,15,25,25,28,16,17,21,20,19,27,21,20,21,19,18,21,20);
		wait for 10 ns;
		t_blur_matrix_int <= (137,136,136,136,132,136,147,148,137,134,133,134,135,141,146,147,135,132,135,136,137,145,146,146,132,137,134,139,144,144,145,142,132,132,135,140,147,149,144,137,135,137,140,142,150,147,138,131,136,137,146,148,147,144,134,128,137,141,146,151,146,139,130,120);
		wait for 10 ns;
		t_blur_matrix_int <= (149,137,129,125,119,119,116,120,146,133,127,116,115,112,110,112,138,127,120,114,108,105,109,107,134,128,115,107,96,93,101,108,128,119,108,100,87,91,95,112,121,114,98,86,83,82,101,118,121,104,87,73,68,79,96,113,112,94,74,64,64,85,99,117);
		wait for 10 ns;
		t_blur_matrix_int <= (119,128,139,137,137,134,134,134,117,129,138,142,137,137,136,135,117,130,138,141,141,135,136,137,118,133,138,138,139,137,137,137,122,132,139,141,141,139,139,142,126,134,140,141,142,141,139,138,124,134,140,144,141,141,138,141,126,134,143,143,142,142,142,138);
		wait for 10 ns;
		t_blur_matrix_int <= (138,138,131,125,113,101,93,73,137,138,131,126,115,102,91,69,141,137,134,124,114,102,87,70,141,137,135,126,113,106,86,69,141,139,134,130,116,101,90,66,139,139,133,124,119,104,85,66,135,140,133,131,116,107,90,67,140,139,134,127,117,101,87,70);
		wait for 10 ns;
		t_blur_matrix_int <= (59,54,49,57,59,61,64,66,58,49,54,56,59,61,62,66,55,51,50,53,60,55,67,67,54,45,53,53,57,59,61,64,54,44,46,52,52,58,63,62,52,42,46,49,64,62,64,62,52,50,46,51,58,55,61,67,53,43,47,50,55,54,59,60);
		wait for 10 ns;
		t_blur_matrix_int <= (69,69,69,75,71,69,71,70,70,69,72,69,67,69,70,71,71,70,70,72,69,75,68,67,67,70,64,66,70,70,70,69,65,65,68,64,67,69,69,66,62,65,66,70,63,67,67,62,69,70,65,65,65,67,65,67,61,63,63,62,65,65,66,70);
		wait for 10 ns;
		t_blur_matrix_int <= (66,68,71,70,79,80,77,75,72,69,69,74,75,79,79,81,70,69,74,71,70,77,79,81,74,67,69,72,78,80,87,82,68,74,72,69,72,77,82,77,63,73,74,70,73,79,79,81,68,69,72,73,75,75,77,76,67,67,69,69,73,76,77,80);
		wait for 10 ns;
		t_blur_matrix_int <= (81,85,88,85,90,88,92,90,83,88,87,89,85,86,92,90,83,87,87,89,86,87,90,89,82,87,84,87,89,89,89,90,85,83,85,86,89,85,92,87,83,84,84,85,87,88,86,89,84,84,84,83,87,90,85,87,81,83,80,83,86,89,88,84);
		wait for 10 ns;
		t_blur_matrix_int <= (93,90,91,94,92,93,91,94,95,89,91,91,89,95,93,91,93,94,92,89,89,90,92,94,91,90,95,90,89,89,94,97,91,87,89,88,92,89,97,89,90,89,86,87,86,93,92,91,84,87,92,89,89,87,91,91,88,86,90,86,89,89,89,91);
		wait for 10 ns;
		t_blur_matrix_int <= (90,91,92,93,93,99,91,92,91,102,95,93,96,94,93,94,96,95,92,95,90,96,95,94,96,95,91,91,92,92,94,89,90,89,94,90,95,93,95,92,93,93,90,92,93,93,91,90,90,92,90,94,94,91,84,89,90,90,90,87,89,89,89,118);
		wait for 10 ns;
		t_blur_matrix_int <= (93,89,94,92,94,93,93,97,97,92,92,88,92,94,95,96,94,96,94,92,93,92,92,91,92,89,93,85,91,93,93,94,93,86,89,88,93,93,97,101,88,85,96,90,106,126,125,126,83,101,154,120,128,125,116,110,97,95,97,110,107,103,99,94);
		wait for 10 ns;
		t_blur_matrix_int <= (98,95,92,95,93,95,88,90,102,92,93,93,92,89,90,90,94,94,91,91,91,89,103,115,91,89,89,97,95,102,120,126,112,111,106,96,99,115,128,117,113,103,87,89,105,104,109,113,98,98,91,91,95,99,108,107,97,92,91,92,95,104,110,109);
		wait for 10 ns;
		t_blur_matrix_int <= (93,92,104,106,113,113,126,125,103,119,122,129,125,130,130,131,118,124,125,134,121,115,124,122,113,122,127,132,122,117,115,129,122,120,122,117,121,122,130,130,113,120,115,114,117,130,124,131,111,102,107,105,122,112,117,129,108,103,101,104,117,104,113,120);
		wait for 10 ns;
		t_blur_matrix_int <= (124,123,126,136,149,145,148,165,128,127,144,160,143,152,152,157,123,138,148,156,156,152,156,163,130,129,140,148,140,147,151,155,120,130,129,133,144,136,146,147,120,129,134,141,136,147,152,153,123,132,128,131,132,148,143,146,126,136,131,135,141,149,141,142);
		wait for 10 ns;
		t_blur_matrix_int <= (161,163,158,173,164,179,168,176,166,172,168,162,165,169,167,165,170,167,165,164,173,153,156,159,161,163,174,166,163,160,162,159,148,159,162,168,162,167,161,170,148,149,163,155,151,168,166,154,158,154,148,151,161,164,172,163,152,148,159,155,166,172,156,178);
		wait for 10 ns;
		t_blur_matrix_int <= (177,163,166,151,118,96,86,85,164,175,182,180,179,164,148,112,170,167,169,179,173,185,183,178,164,175,167,171,177,179,176,188,157,170,173,168,172,180,179,179,172,168,171,184,174,179,185,182,158,180,173,172,183,177,176,182,178,172,177,175,164,177,184,174);
		wait for 10 ns;
		t_blur_matrix_int <= (85,87,86,93,90,89,92,93,91,86,78,85,85,90,88,88,165,132,100,80,82,82,89,88,183,184,170,124,84,80,84,85,186,193,186,182,158,105,80,79,181,186,188,186,185,180,125,84,186,185,180,186,192,189,186,156,176,187,185,184,188,193,193,186);
		wait for 10 ns;
		t_blur_matrix_int <= (95,101,99,97,100,98,95,91,94,96,99,97,95,94,95,91,91,92,96,91,90,92,94,92,82,92,92,93,90,94,92,97,85,88,94,90,96,95,94,92,76,87,90,87,89,94,91,87,104,80,88,79,82,82,87,88,176,129,88,77,79,80,85,84);
		wait for 10 ns;
		t_blur_matrix_int <= (98,89,94,93,91,96,91,91,93,91,90,92,91,91,91,91,92,92,91,95,87,88,89,93,91,91,90,93,90,90,90,87,89,90,89,93,89,90,86,88,86,87,92,87,87,89,87,86,88,87,88,87,86,84,88,88,84,84,90,85,87,84,86,86);
		wait for 10 ns;
		t_blur_matrix_int <= (93,89,88,84,88,85,78,78,88,85,84,85,83,86,82,77,87,83,86,84,82,83,83,77,88,84,87,83,82,80,81,78,87,85,82,83,77,82,81,78,83,82,82,79,78,76,79,74,86,84,80,80,79,80,78,77,86,84,84,80,77,79,74,74);
		wait for 10 ns;
		t_blur_matrix_int <= (78,79,76,73,75,79,86,92,79,76,76,75,74,80,85,95,80,82,74,71,72,78,88,99,80,80,74,73,80,77,89,95,81,75,78,73,79,78,90,93,76,70,70,72,78,79,82,92,76,75,68,68,74,78,81,95,75,70,69,64,74,75,85,93);
		wait for 10 ns;
		t_blur_matrix_int <= (100,107,113,115,113,116,120,115,102,109,114,116,115,114,116,117,102,110,110,121,114,115,113,116,104,107,114,115,116,114,115,115,106,112,109,114,119,116,114,115,103,108,114,118,116,117,116,115,100,112,114,116,116,117,116,114,104,107,111,118,118,116,115,115);
		wait for 10 ns;
		t_blur_matrix_int <= (122,122,125,127,127,128,128,128,118,121,122,123,128,126,127,128,118,119,119,123,122,130,125,126,118,118,119,121,124,126,125,127,116,118,121,118,124,122,123,123,116,115,118,121,118,120,124,125,111,119,118,117,114,117,125,125,115,116,119,118,119,117,118,122);
		wait for 10 ns;
		t_blur_matrix_int <= (122,125,125,126,124,127,128,127,125,127,127,127,127,123,126,123,128,122,123,123,126,123,123,124,126,124,121,123,126,123,121,118,124,124,121,119,120,119,119,118,125,123,122,117,119,117,118,119,121,124,125,121,116,112,116,113,119,121,124,125,119,117,114,109);
		wait for 10 ns;
		t_blur_matrix_int <= (126,127,123,123,122,124,121,120,126,129,122,124,123,117,117,119,122,123,121,122,116,117,115,114,117,122,117,119,115,116,113,112,116,120,118,115,116,114,113,116,114,114,119,116,115,116,112,111,111,115,113,116,117,117,113,113,109,113,114,115,117,117,113,115);
		wait for 10 ns;
		t_blur_matrix_int <= (118,115,118,115,117,114,112,114,116,113,113,115,111,111,111,112,116,110,111,112,111,109,111,112,118,115,110,110,111,108,109,112,112,111,113,106,110,107,107,111,112,111,111,111,110,112,108,108,110,112,111,113,111,108,112,111,112,114,116,111,111,111,111,112);
		wait for 10 ns;
		t_blur_matrix_int <= (114,113,114,111,117,119,161,191,111,112,111,109,111,118,131,176,113,115,115,111,112,113,116,150,114,111,112,109,111,114,107,117,110,112,112,112,111,113,107,107,108,108,112,109,111,114,109,108,109,111,112,113,112,114,112,108,111,112,114,113,114,113,108,111);
		wait for 10 ns;
		t_blur_matrix_int <= (205,212,215,219,218,219,208,179,197,208,213,218,221,223,216,201,187,202,210,215,220,222,223,213,171,196,208,216,219,220,223,221,136,182,203,214,218,220,222,224,113,158,196,207,214,219,223,223,105,125,176,196,210,217,221,224,112,115,149,188,207,215,222,226);
		wait for 10 ns;
		t_blur_matrix_int <= (119,79,74,84,85,95,82,63,161,98,80,88,93,86,61,27,193,141,90,89,88,71,29,19,210,183,117,91,67,33,21,15,221,205,158,77,35,16,18,18,224,216,189,71,17,17,14,16,228,222,188,47,9,18,14,16,225,212,124,14,15,17,18,18);
		wait for 10 ns;
		t_blur_matrix_int <= (28,13,19,17,17,21,18,22,17,16,15,18,17,17,20,20,14,13,20,17,19,22,18,22,17,20,24,24,23,27,25,30,15,16,20,21,30,31,28,24,20,20,22,18,24,29,23,25,20,23,21,22,29,28,27,24,18,19,21,26,29,27,25,28);
		wait for 10 ns;
		t_blur_matrix_int <= (25,34,25,36,36,34,34,30,30,25,27,26,26,29,28,28,29,30,25,25,27,23,25,26,29,31,26,26,26,20,18,19,30,25,25,26,23,20,22,28,28,24,29,27,21,27,21,24,28,32,20,19,18,21,25,35,27,21,19,19,16,24,32,23);
		wait for 10 ns;
		t_blur_matrix_int <= (24,15,16,17,22,19,22,21,22,16,17,14,17,18,17,20,22,20,25,23,22,17,17,16,28,29,22,20,21,19,18,22,31,24,19,21,17,19,24,18,25,20,22,24,23,18,18,22,26,23,17,28,24,18,26,24,19,20,19,20,20,23,32,29);
		wait for 10 ns;
		t_blur_matrix_int <= (141,147,155,149,144,131,127,117,146,152,154,148,137,131,119,113,147,149,150,141,133,125,116,99,150,147,145,139,132,120,108,89,147,148,145,133,126,114,98,84,149,146,136,130,119,108,85,68,144,140,133,125,113,96,77,53,140,134,127,118,104,86,63,45);
		wait for 10 ns;
		t_blur_matrix_int <= (105,81,65,50,56,81,98,115,95,74,58,42,62,80,101,115,85,59,40,42,59,81,98,111,70,44,42,47,63,82,98,111,58,46,40,51,65,79,98,111,48,44,42,51,65,85,99,109,57,50,43,52,67,86,99,112,50,54,49,47,64,83,98,113);
		wait for 10 ns;
		t_blur_matrix_int <= (127,134,141,142,143,142,141,140,126,139,142,143,142,143,144,136,125,139,140,145,142,137,140,138,121,136,142,145,144,137,141,141,123,135,143,145,145,142,142,139,127,137,142,145,143,142,141,138,123,137,142,143,142,143,142,138,124,134,141,144,146,145,145,140);
		wait for 10 ns;
		t_blur_matrix_int <= (140,138,138,124,117,102,86,67,137,137,134,121,114,102,86,70,138,137,131,124,109,98,84,66,139,139,130,122,108,101,84,69,137,134,132,122,111,102,84,66,139,137,131,119,114,98,86,67,136,134,132,123,114,97,86,62,137,134,133,126,113,102,83,68);
		wait for 10 ns;
		t_blur_matrix_int <= (51,43,45,50,48,51,57,63,50,44,41,45,52,56,63,59,52,41,40,49,54,56,60,63,47,40,40,50,56,52,59,64,44,44,38,49,53,58,61,63,43,42,42,50,54,57,63,60,45,41,42,49,51,51,63,62,50,39,46,49,57,53,63,69);
		wait for 10 ns;
		t_blur_matrix_int <= (63,63,60,67,65,67,66,66,58,62,63,61,63,67,66,67,60,66,68,64,65,67,65,67,70,72,70,72,66,70,68,65,67,68,66,74,67,67,60,66,66,64,68,71,66,72,66,68,71,63,62,63,65,68,66,67,72,66,64,68,68,65,68,65);
		wait for 10 ns;
		t_blur_matrix_int <= (70,69,69,71,72,78,70,79,68,68,71,66,71,69,68,78,71,67,68,69,73,75,74,78,69,67,72,67,74,74,73,78,64,69,62,70,72,75,76,75,65,65,68,68,72,72,77,75,69,69,67,70,71,74,75,78,69,67,68,71,70,73,78,81);
		wait for 10 ns;
		t_blur_matrix_int <= (82,82,84,82,85,84,84,82,79,80,80,81,85,80,81,83,79,79,78,79,80,83,84,83,82,84,74,77,83,82,85,85,80,77,83,83,84,81,82,82,81,79,80,80,77,80,83,87,77,78,82,84,80,81,82,90,83,85,84,78,79,79,85,80);
		wait for 10 ns;
		t_blur_matrix_int <= (90,87,91,89,86,87,94,90,96,90,88,90,91,89,90,86,86,86,86,85,89,89,86,93,85,85,83,85,86,87,91,90,87,85,84,85,87,85,88,87,86,83,85,85,88,87,89,88,84,82,88,83,88,87,82,87,88,83,86,86,88,84,87,85);
		wait for 10 ns;
		t_blur_matrix_int <= (90,86,90,86,89,86,102,154,89,90,91,88,79,88,156,110,89,90,89,87,92,87,116,82,89,86,90,88,90,112,79,77,89,84,86,83,112,98,77,80,89,88,86,101,166,81,77,84,93,87,84,119,110,77,81,78,86,86,91,119,85,83,76,73);
		wait for 10 ns;
		t_blur_matrix_int <= (77,86,94,91,95,95,89,92,58,79,92,90,96,88,93,87,73,79,84,85,94,86,87,95,82,75,85,87,86,86,90,89,83,84,82,80,76,82,84,86,80,78,76,75,79,83,86,89,73,74,74,80,80,87,89,85,70,75,74,84,87,88,83,85);
		wait for 10 ns;
		t_blur_matrix_int <= (92,90,97,92,98,109,110,107,96,91,91,87,97,107,102,107,101,91,87,93,99,101,104,107,95,92,92,91,101,107,110,107,94,92,97,94,96,105,93,103,96,103,91,96,103,96,92,103,93,86,99,98,92,94,102,108,79,99,90,99,88,97,104,100);
		wait for 10 ns;
		t_blur_matrix_int <= (105,99,105,111,116,113,111,117,100,103,104,109,108,107,116,109,103,101,101,106,111,113,106,107,101,106,107,111,111,106,97,107,109,105,108,109,110,99,102,114,107,105,111,109,106,108,115,108,100,104,98,109,113,110,112,107,100,96,103,108,105,109,107,105);
		wait for 10 ns;
		t_blur_matrix_int <= (124,124,116,133,132,146,133,136,119,114,122,133,130,131,140,137,112,119,120,118,128,134,136,146,115,106,106,122,120,134,138,146,110,124,114,124,124,119,140,133,112,107,120,111,124,131,122,141,108,115,100,120,126,123,127,127,114,114,115,122,122,121,126,124);
		wait for 10 ns;
		t_blur_matrix_int <= (150,141,166,155,154,166,173,177,164,157,156,162,163,165,176,174,147,164,161,159,163,163,165,171,150,154,163,161,153,172,164,159,149,151,144,162,152,156,173,176,134,150,145,141,159,170,160,167,145,129,153,164,153,166,172,169,139,149,149,151,172,169,167,180);
		wait for 10 ns;
		t_blur_matrix_int <= (179,176,165,175,177,178,181,181,163,180,180,168,177,184,174,169,173,170,176,175,174,171,185,180,168,175,162,167,184,182,177,184,169,169,179,183,176,183,184,181,176,167,174,178,186,179,178,186,169,180,177,168,178,184,180,175,181,171,167,183,176,167,183,186);
		wait for 10 ns;
		t_blur_matrix_int <= (176,173,185,187,186,184,187,190,180,185,180,186,191,187,187,186,175,179,184,184,184,188,192,188,186,176,181,190,188,186,188,191,180,188,183,185,186,191,186,187,183,180,186,192,183,186,188,186,183,184,187,184,187,188,184,182,182,174,189,188,179,182,182,173);
		wait for 10 ns;
		t_blur_matrix_int <= (189,183,149,99,75,77,77,78,187,184,187,173,116,76,69,73,182,189,190,193,189,150,87,68,190,186,189,195,194,193,160,89,184,193,191,193,194,194,196,165,187,187,189,189,182,179,189,198,186,184,171,176,188,198,206,212,173,184,195,205,206,207,211,211);
		wait for 10 ns;
		t_blur_matrix_int <= (83,89,84,84,83,84,83,82,79,86,79,79,82,82,82,84,77,73,71,72,76,80,80,80,66,65,72,71,74,73,76,79,99,60,65,62,64,67,72,76,176,127,114,82,59,64,66,70,217,218,215,189,95,54,58,69,213,221,224,224,179,67,52,55);
		wait for 10 ns;
		t_blur_matrix_int <= (83,83,83,82,77,79,76,80,81,82,80,76,78,73,76,75,80,79,79,78,76,80,78,72,82,78,79,78,77,76,75,74,81,75,81,75,73,71,75,76,78,75,78,74,73,75,70,70,77,72,74,76,71,68,71,71,68,70,75,72,68,67,67,69);
		wait for 10 ns;
		t_blur_matrix_int <= (70,75,70,68,69,75,83,95,74,71,68,66,69,79,87,93,73,73,72,69,70,78,80,96,72,75,72,65,70,74,82,89,79,72,69,66,69,73,83,94,73,67,67,65,66,76,78,94,73,69,71,65,69,75,83,97,71,69,69,62,71,73,78,94);
		wait for 10 ns;
		t_blur_matrix_int <= (102,108,115,118,121,117,117,115,105,109,117,119,120,121,119,115,105,113,117,122,123,121,120,119,105,109,119,123,120,123,120,123,105,113,117,125,122,124,125,120,110,118,122,124,125,128,128,125,109,114,123,125,126,128,128,125,108,116,119,123,129,125,128,123);
		wait for 10 ns;
		t_blur_matrix_int <= (116,112,116,114,116,115,117,116,116,115,114,116,113,113,111,111,117,114,115,114,109,116,109,111,120,120,114,109,106,108,106,106,121,116,114,109,102,102,102,99,119,119,120,110,101,97,91,93,122,124,120,110,100,92,86,79,122,123,124,114,102,87,80,68);
		wait for 10 ns;
		t_blur_matrix_int <= (117,124,123,121,120,112,111,110,117,116,120,123,123,113,111,108,108,111,114,123,122,114,116,112,103,106,110,119,120,118,115,112,98,98,103,111,120,121,118,115,89,92,97,110,115,121,118,115,84,83,95,100,112,116,120,117,74,73,83,93,106,111,119,119);
		wait for 10 ns;
		t_blur_matrix_int <= (110,112,109,112,112,118,112,110,111,109,111,112,116,116,116,112,108,112,114,114,115,117,116,111,112,112,113,111,114,116,115,112,110,110,112,113,116,116,114,112,112,110,113,116,116,120,119,108,112,114,115,114,120,117,116,110,115,114,113,114,114,116,115,112);
		wait for 10 ns;
		t_blur_matrix_int <= (113,114,114,111,111,107,112,109,110,114,111,112,112,111,113,111,113,111,112,112,111,111,112,112,111,112,111,111,111,110,115,112,111,112,112,110,111,114,113,115,110,111,109,111,112,111,114,115,110,111,112,111,112,112,114,113,110,114,110,113,110,112,112,112);
		wait for 10 ns;
		t_blur_matrix_int <= (107,112,117,114,115,117,113,112,111,111,115,116,112,115,116,113,112,114,112,114,111,114,116,117,114,116,110,115,115,116,114,118,114,115,113,118,112,116,120,121,115,113,116,122,117,118,120,119,113,115,116,113,112,117,119,119,111,111,115,114,117,119,118,122);
		wait for 10 ns;
		t_blur_matrix_int <= (113,111,121,164,201,215,223,224,117,114,116,131,190,209,220,208,117,120,121,119,161,200,204,167,116,122,123,123,145,179,143,59,120,119,126,126,131,111,50,22,120,123,127,127,107,56,23,20,122,128,129,119,75,23,19,20,125,127,123,86,38,24,17,21);
		wait for 10 ns;
		t_blur_matrix_int <= (212,165,40,12,17,12,14,17,170,66,16,16,18,19,19,17,72,16,16,19,21,16,18,18,20,20,21,19,19,19,20,23,20,19,22,17,21,23,21,25,18,17,20,15,14,18,25,30,19,17,18,17,18,27,23,27,21,11,25,16,19,24,24,23);
		wait for 10 ns;
		t_blur_matrix_int <= (24,21,23,31,26,24,28,29,23,20,29,32,26,31,30,28,21,27,21,21,29,28,28,22,22,21,24,25,28,26,23,19,27,25,25,26,23,25,18,16,32,25,23,21,18,19,12,18,29,29,25,18,16,20,22,29,26,22,16,18,16,22,26,31);
		wait for 10 ns;
		t_blur_matrix_int <= (24,17,18,17,20,25,25,26,27,14,18,23,23,29,22,16,20,22,22,26,28,22,20,20,24,31,29,28,26,27,19,24,24,35,25,23,27,22,20,28,26,27,31,29,20,28,26,30,31,29,24,25,23,23,27,32,25,29,24,23,22,26,35,45);
		wait for 10 ns;
		t_blur_matrix_int <= (22,17,17,19,22,29,22,16,20,19,24,26,28,27,15,7,19,17,31,34,33,18,9,6,23,24,40,45,29,11,5,15,30,40,45,30,18,9,13,70,36,43,33,16,7,13,58,116,50,37,17,14,13,48,105,137,55,31,14,19,40,88,126,144);
		wait for 10 ns;
		t_blur_matrix_int <= (133,133,121,109,93,77,58,45,135,127,116,99,81,64,46,48,124,121,107,91,69,52,47,53,117,113,96,75,56,44,54,53,113,103,84,62,49,49,55,56,101,93,70,54,49,54,55,53,90,81,60,49,54,55,63,55,82,67,50,50,53,61,63,57);
		wait for 10 ns;
		t_blur_matrix_int <= (49,52,52,50,69,87,100,115,53,50,49,51,67,84,100,113,52,52,54,56,67,83,97,113,58,58,48,59,66,84,100,111,56,52,48,56,69,84,101,115,58,54,55,52,69,81,96,113,58,53,56,54,62,84,94,114,56,56,49,52,64,81,99,113);
		wait for 10 ns;
		t_blur_matrix_int <= (124,135,138,143,144,142,144,141,124,133,139,146,143,144,144,142,124,132,141,145,146,145,143,142,124,136,141,143,144,143,140,141,123,134,140,143,143,141,140,142,121,129,138,140,145,142,141,140,122,132,138,139,143,145,139,138,120,128,137,139,145,143,141,143);
		wait for 10 ns;
		t_blur_matrix_int <= (140,139,132,123,112,96,82,63,141,133,131,120,109,98,79,62,140,135,127,121,109,96,76,76,142,139,130,122,109,98,83,69,145,138,129,121,110,97,81,66,138,140,130,121,110,95,78,69,139,136,133,122,108,94,82,62,140,135,131,124,110,96,78,64);
		wait for 10 ns;
		t_blur_matrix_int <= (53,43,38,49,51,56,59,62,48,41,42,50,55,58,61,62,53,43,43,50,53,56,63,63,53,44,50,51,58,56,57,61,53,44,39,49,50,58,60,64,49,40,45,52,58,58,62,65,54,43,43,56,54,61,64,65,50,42,49,52,59,66,65,66);
		wait for 10 ns;
		t_blur_matrix_int <= (62,63,64,62,69,68,64,69,60,70,68,67,67,67,67,64,63,66,63,66,67,64,76,71,64,64,67,65,66,69,74,67,59,61,63,70,69,70,71,70,61,63,68,71,67,71,71,66,65,59,62,68,65,63,67,63,70,65,65,66,64,67,67,67);
		wait for 10 ns;
		t_blur_matrix_int <= (69,68,67,69,73,76,78,76,65,69,72,72,72,75,76,80,67,69,65,71,66,73,78,79,66,65,67,69,72,74,75,75,69,66,68,69,75,76,74,75,68,66,66,73,72,73,73,75,64,65,69,72,72,70,72,81,69,67,66,73,72,71,75,77);
		wait for 10 ns;
		t_blur_matrix_int <= (77,80,82,80,80,86,87,90,79,79,82,81,80,82,83,88,80,82,81,82,81,85,82,88,77,81,80,79,81,81,82,85,79,79,82,82,82,81,86,85,80,80,83,83,80,83,88,90,79,79,84,82,82,84,85,85,81,79,82,85,80,83,83,83);
		wait for 10 ns;
		t_blur_matrix_int <= (87,86,91,86,91,87,82,84,85,83,90,87,88,84,89,86,84,87,88,86,90,86,93,89,85,84,85,86,90,90,92,89,86,86,88,86,89,88,93,95,88,87,80,91,85,87,94,88,83,91,86,86,89,90,91,77,85,85,90,90,90,93,84,84);
		wait for 10 ns;
		t_blur_matrix_int <= (90,89,103,91,80,76,71,77,90,92,92,81,74,75,77,76,91,96,81,72,76,73,75,76,93,86,77,70,71,71,80,81,81,79,74,74,76,72,81,83,74,76,70,74,79,76,80,81,73,74,75,77,80,80,78,77,74,72,77,83,81,76,85,81);
		wait for 10 ns;
		t_blur_matrix_int <= (74,78,78,83,92,81,81,87,77,83,85,89,87,80,90,93,78,88,85,84,83,93,90,86,83,88,76,87,95,88,88,90,78,79,85,89,89,84,81,96,77,91,92,81,88,84,89,86,87,88,86,87,86,85,85,78,87,84,86,84,74,82,72,79);
		wait for 10 ns;
		t_blur_matrix_int <= (93,92,91,92,93,94,101,100,88,91,91,90,89,95,84,97,90,90,92,83,95,88,96,95,90,85,90,85,84,94,97,102,84,86,84,84,87,98,94,104,80,81,88,94,89,100,99,87,77,82,94,98,101,97,100,103,84,90,85,101,97,102,97,103);
		wait for 10 ns;
		t_blur_matrix_int <= (98,92,105,100,107,102,114,105,96,102,99,114,98,108,97,111,102,102,105,108,114,105,118,98,107,97,110,116,103,111,107,111,94,107,106,110,105,100,113,102,102,107,118,104,110,116,107,114,103,119,110,115,117,112,120,110,107,105,114,104,116,117,114,119);
		wait for 10 ns;
		t_blur_matrix_int <= (104,104,114,130,107,123,128,138,104,107,114,112,111,105,126,122,111,107,112,114,105,122,116,128,105,113,123,110,117,107,128,133,110,116,108,113,117,127,119,125,112,117,119,113,123,123,123,121,119,119,118,116,113,114,112,118,123,122,111,104,119,108,120,120);
		wait for 10 ns;
		t_blur_matrix_int <= (140,125,159,161,160,174,178,168,136,149,143,152,171,173,162,177,138,134,153,155,155,174,174,168,128,139,145,152,161,171,153,174,134,126,146,148,147,163,169,160,129,140,133,143,164,170,157,165,123,128,145,158,153,160,168,150,123,143,143,145,169,148,141,128);
		wait for 10 ns;
		t_blur_matrix_int <= (166,182,170,167,178,183,175,179,179,168,171,184,172,168,180,185,172,179,186,176,178,180,166,163,170,168,174,183,172,141,149,160,161,179,166,149,148,149,178,191,172,160,132,141,166,183,200,199,138,131,157,189,196,196,191,197,129,163,192,199,198,200,195,186);
		wait for 10 ns;
		t_blur_matrix_int <= (183,186,177,174,176,170,176,190,174,166,161,168,178,193,204,207,156,164,178,196,204,206,202,204,183,200,203,211,202,200,195,197,205,205,204,202,200,198,193,197,203,202,197,195,195,197,201,192,191,193,198,203,207,199,195,195,195,197,203,203,196,199,191,194);
		wait for 10 ns;
		t_blur_matrix_int <= (203,207,204,204,211,206,206,209,208,201,204,202,203,208,202,205,203,202,200,205,201,203,205,198,200,204,203,198,199,198,203,207,202,197,200,200,195,201,198,200,199,201,200,199,198,195,198,198,191,195,195,193,193,195,199,206,187,182,188,198,194,202,209,212);
		wait for 10 ns;
		t_blur_matrix_int <= (211,214,222,225,218,126,49,51,210,208,218,222,222,196,93,48,202,207,210,219,218,224,179,67,197,202,210,212,219,217,216,146,207,197,202,204,208,223,217,212,199,205,208,209,211,221,224,216,205,209,209,211,212,219,224,220,206,201,204,200,204,209,211,222);
		wait for 10 ns;
		t_blur_matrix_int <= (62,65,70,68,72,68,69,70,55,61,69,65,69,67,68,65,49,54,59,62,61,67,63,64,57,45,50,58,62,67,65,64,136,50,47,49,57,60,66,63,198,91,46,48,52,55,55,63,218,178,65,44,50,47,54,56,218,219,133,64,48,44,51,51);
		wait for 10 ns;
		t_blur_matrix_int <= (65,67,67,64,68,78,80,96,70,68,66,61,66,75,79,96,69,63,64,64,62,74,81,93,68,64,63,57,65,72,79,91,65,63,64,62,63,71,80,90,67,62,64,59,64,69,82,92,56,58,59,59,64,71,81,92,55,56,55,54,63,72,81,93);
		wait for 10 ns;
		t_blur_matrix_int <= (102,114,119,123,127,124,127,125,105,112,117,122,126,122,126,124,101,110,119,129,126,123,123,122,100,112,121,126,126,123,122,124,104,111,121,126,124,125,126,122,99,111,119,126,127,128,126,123,105,113,123,125,127,124,126,124,105,112,120,126,126,124,125,122);
		wait for 10 ns;
		t_blur_matrix_int <= (123,124,124,113,103,90,74,62,122,124,122,115,108,96,78,54,125,123,120,113,107,95,78,57,124,123,122,112,106,99,81,55,123,120,121,117,107,96,85,64,123,121,123,120,112,100,86,65,125,124,123,115,111,103,89,66,125,126,123,118,112,98,85,59);
		wait for 10 ns;
		t_blur_matrix_int <= (59,59,73,85,98,106,115,120,49,49,53,73,89,105,109,114,37,33,40,64,83,98,103,112,27,23,25,52,75,88,102,108,35,18,22,35,59,80,91,104,35,13,16,23,48,71,80,95,35,16,15,24,42,68,75,88,37,13,14,20,36,60,71,86);
		wait for 10 ns;
		t_blur_matrix_int <= (117,114,111,112,110,116,113,112,118,115,115,110,115,116,114,112,118,116,116,110,113,118,115,114,117,118,118,113,111,111,114,115,112,117,122,117,111,112,110,116,106,116,118,119,113,111,113,111,102,110,115,118,115,111,115,112,99,105,111,118,117,117,113,112);
		wait for 10 ns;
		t_blur_matrix_int <= (112,110,113,111,112,117,113,116,111,110,114,112,111,112,113,117,111,113,114,110,109,113,115,111,109,109,114,112,112,110,113,112,113,112,112,112,111,114,112,115,112,109,112,109,115,110,112,114,110,112,111,109,114,110,114,114,107,114,107,112,112,111,112,112);
		wait for 10 ns;
		t_blur_matrix_int <= (115,114,114,114,115,119,115,121,112,114,114,114,118,116,118,126,113,111,115,116,120,119,120,126,110,111,113,110,111,121,125,123,109,114,111,114,117,122,125,108,111,117,118,117,120,126,114,66,113,113,117,117,125,127,90,31,113,114,115,119,123,108,55,17);
		wait for 10 ns;
		t_blur_matrix_int <= (127,122,95,46,16,26,18,23,129,108,61,21,18,17,11,13,118,77,29,16,16,12,12,16,99,36,16,10,15,13,13,14,52,20,17,16,18,17,17,22,22,20,55,47,30,17,18,28,20,18,19,22,17,16,20,22,13,12,20,17,19,23,26,26);
		wait for 10 ns;
		t_blur_matrix_int <= (17,19,24,21,23,31,21,28,14,16,20,23,24,29,27,24,20,21,27,27,28,23,27,23,19,25,25,27,27,27,28,25,30,30,28,29,27,28,23,22,30,25,25,27,29,25,22,23,25,25,21,26,24,22,20,20,27,25,31,27,18,18,12,18);
		wait for 10 ns;
		t_blur_matrix_int <= (26,23,25,18,16,29,27,31,23,19,18,16,21,29,29,24,23,18,19,24,25,27,25,19,18,12,25,26,28,25,20,20,21,18,33,33,25,19,18,20,20,26,29,30,22,24,23,23,24,32,34,20,24,29,24,25,30,29,30,18,23,24,26,23);
		wait for 10 ns;
		t_blur_matrix_int <= (21,22,24,18,21,31,45,58,20,23,24,21,29,40,44,48,20,21,27,26,34,49,54,39,22,28,47,50,39,53,48,41,25,34,39,39,45,55,47,51,24,35,36,43,51,49,58,75,24,34,42,45,56,57,74,97,30,31,38,52,56,79,98,118);
		wait for 10 ns;
		t_blur_matrix_int <= (53,29,18,41,87,119,131,146,43,24,38,81,113,125,134,137,36,49,79,110,125,125,125,133,50,76,106,124,130,122,122,125,80,105,122,129,129,119,114,116,102,117,124,128,130,113,109,129,116,121,126,128,124,111,126,139,126,127,122,124,112,122,139,144);
		wait for 10 ns;
		t_blur_matrix_int <= (67,57,50,53,53,56,58,59,59,50,53,54,55,59,62,58,57,52,55,59,54,57,56,56,60,55,56,60,61,59,58,61,52,55,58,59,59,60,60,62,53,52,59,61,60,58,61,64,58,57,57,62,59,62,57,55,62,60,57,59,60,56,58,62);
		wait for 10 ns;
		t_blur_matrix_int <= (57,54,49,56,61,80,98,109,60,56,51,52,67,79,94,107,60,56,52,54,62,78,92,112,58,58,54,56,65,77,98,111,59,59,54,61,65,84,97,111,61,58,57,59,71,82,99,108,58,57,54,52,67,83,95,110,60,54,55,54,65,78,96,112);
		wait for 10 ns;
		t_blur_matrix_int <= (120,130,135,140,141,142,143,140,119,130,135,138,142,139,141,139,117,131,134,139,141,140,140,141,117,129,136,140,141,142,146,141,116,130,133,136,143,140,140,138,118,130,133,138,137,135,138,142,121,130,135,138,142,138,139,137,119,129,133,137,139,141,141,135);
		wait for 10 ns;
		t_blur_matrix_int <= (138,138,130,125,109,101,82,76,136,134,133,120,106,93,83,67,140,139,132,122,111,97,82,66,140,136,130,122,111,94,83,70,137,135,131,121,111,97,82,65,133,137,131,123,112,101,81,67,139,139,134,124,112,98,82,69,135,138,136,124,114,101,86,69);
		wait for 10 ns;
		t_blur_matrix_int <= (50,42,52,54,59,59,66,63,56,42,43,42,56,59,63,63,52,43,44,46,56,56,62,63,61,41,40,49,50,58,61,60,59,41,44,47,55,60,64,62,54,44,43,47,53,58,60,61,61,43,45,50,53,56,60,60,53,43,45,49,54,51,59,60);
		wait for 10 ns;
		t_blur_matrix_int <= (68,69,63,65,64,64,66,68,65,68,66,68,64,65,64,66,65,69,67,66,67,70,63,71,66,63,64,66,65,69,67,68,65,61,62,69,72,65,63,66,59,62,63,66,69,66,67,63,65,68,66,65,67,67,70,66,63,65,65,66,69,68,69,69);
		wait for 10 ns;
		t_blur_matrix_int <= (65,71,69,70,70,70,74,79,67,65,70,69,75,72,74,77,65,72,72,68,70,72,77,74,70,69,65,68,69,74,76,76,67,68,66,68,69,73,75,73,62,67,68,69,69,71,75,76,64,65,69,68,69,72,73,78,67,68,68,69,76,77,78,74);
		wait for 10 ns;
		t_blur_matrix_int <= (78,81,88,85,82,83,80,86,79,83,83,82,83,79,84,85,77,80,84,82,83,86,83,84,78,83,85,85,88,84,86,84,77,80,80,85,85,87,85,81,78,76,80,84,81,80,80,78,82,80,82,82,79,83,79,79,80,76,78,81,84,80,73,75);
		wait for 10 ns;
		t_blur_matrix_int <= (86,86,87,90,97,89,88,81,88,86,88,93,102,80,79,75,88,83,86,104,95,72,71,73,85,86,99,100,82,75,80,69,79,91,138,83,70,65,68,70,77,132,144,77,65,68,73,68,84,167,131,68,60,67,75,72,108,187,116,65,66,68,71,75);
		wait for 10 ns;
		t_blur_matrix_int <= (79,85,72,82,77,79,82,83,81,84,79,80,76,82,81,83,75,84,78,78,77,77,79,81,76,79,83,78,83,77,81,82,70,77,81,85,82,75,82,79,74,78,77,81,80,77,79,80,78,81,76,81,77,79,76,80,75,74,75,79,74,80,83,79);
		wait for 10 ns;
		t_blur_matrix_int <= (88,84,82,79,81,87,86,90,86,84,80,87,87,92,87,87,84,86,78,88,87,86,87,88,78,81,84,85,80,88,88,94,84,83,81,82,89,84,87,95,80,78,79,80,87,91,94,89,76,84,85,88,86,95,94,88,89,91,86,88,90,89,98,94);
		wait for 10 ns;
		t_blur_matrix_int <= (88,91,96,91,107,94,104,101,90,90,101,102,97,106,96,107,95,100,97,103,97,96,110,102,102,103,103,93,108,111,107,119,104,97,102,114,104,117,118,110,92,109,105,96,116,114,115,114,98,92,107,105,111,122,103,96,97,103,110,111,118,97,104,105);
		wait for 10 ns;
		t_blur_matrix_int <= (111,108,98,113,111,116,115,120,116,106,116,102,110,115,105,117,111,111,102,109,112,117,112,111,115,104,123,106,109,109,108,111,114,108,109,119,113,109,116,102,91,110,113,111,121,108,113,113,108,107,105,116,105,111,108,99,105,105,115,107,113,108,100,102);
		wait for 10 ns;
		t_blur_matrix_int <= (122,108,113,114,110,114,116,120,110,115,109,104,114,110,124,119,108,109,105,106,109,114,109,119,101,108,103,98,112,111,117,110,109,107,108,104,109,113,107,101,99,105,92,99,107,96,97,100,108,94,96,94,97,91,116,156,96,100,81,80,85,131,158,153);
		wait for 10 ns;
		t_blur_matrix_int <= (130,128,146,158,145,120,115,148,117,140,150,137,111,110,166,178,126,139,129,105,129,177,190,180,106,114,109,145,178,186,188,189,105,124,154,166,181,182,190,190,150,177,167,162,171,187,188,188,159,185,172,174,177,178,178,182,175,175,192,176,179,167,173,175);
		wait for 10 ns;
		t_blur_matrix_int <= (172,195,193,194,193,194,194,194,187,185,195,193,185,197,200,200,180,185,182,197,191,187,196,192,182,186,189,178,185,186,182,185,190,175,184,183,176,183,184,179,179,185,177,184,181,175,186,179,177,182,185,173,184,178,168,175,184,185,179,174,159,182,183,186);
		wait for 10 ns;
		t_blur_matrix_int <= (195,202,189,195,192,185,187,188,189,185,197,190,180,190,184,195,192,185,186,193,187,198,181,187,187,187,193,192,188,180,189,195,186,186,179,182,192,197,196,190,166,178,183,192,195,196,195,197,179,187,192,188,194,196,196,198,189,183,187,193,187,194,197,197);
		wait for 10 ns;
		t_blur_matrix_int <= (200,194,195,203,195,193,197,192,201,197,189,190,188,193,195,196,187,191,197,196,196,197,199,197,200,189,195,205,199,200,197,200,199,201,189,198,201,201,200,198,186,199,200,192,198,194,199,195,200,190,205,193,189,201,200,198,198,191,193,201,193,195,197,197);
		wait for 10 ns;
		t_blur_matrix_int <= (194,196,198,200,201,207,208,209,193,201,203,203,206,205,205,206,197,201,202,203,202,206,203,205,202,201,199,201,202,203,204,198,199,202,196,197,202,203,203,199,202,205,200,201,201,202,199,201,199,200,199,199,199,196,196,195,197,196,193,191,194,201,199,201);
		wait for 10 ns;
		t_blur_matrix_int <= (211,216,206,159,95,62,43,46,209,214,217,221,206,132,51,44,209,210,213,219,221,214,139,71,207,207,206,205,211,223,213,124,206,210,208,209,207,214,216,206,197,209,209,209,211,217,210,215,195,202,207,211,209,219,216,221,198,203,206,209,210,210,220,222);
		wait for 10 ns;
		t_blur_matrix_int <= (48,50,57,52,58,67,81,93,39,49,50,52,56,66,78,92,35,41,46,48,55,65,78,88,38,32,39,45,54,63,77,95,85,24,33,40,53,61,78,90,174,41,32,35,46,58,72,90,209,101,59,31,41,55,71,85,225,196,87,27,39,51,71,90);
		wait for 10 ns;
		t_blur_matrix_int <= (103,110,119,126,125,125,125,121,104,112,118,127,125,125,128,126,104,114,121,126,127,123,126,123,102,111,121,127,124,125,125,122,99,110,120,121,125,123,121,125,99,110,118,124,124,124,125,126,98,110,118,122,125,124,127,125,100,109,116,122,122,122,126,125);
		wait for 10 ns;
		t_blur_matrix_int <= (123,126,121,118,112,100,89,60,124,122,125,121,114,99,86,60,120,126,126,131,108,100,81,65,123,122,128,120,108,99,82,64,122,123,125,119,109,100,84,67,123,125,122,118,111,98,88,69,122,125,122,119,106,99,83,66,126,124,124,120,110,98,83,67);
		wait for 10 ns;
		t_blur_matrix_int <= (34,15,24,25,32,50,66,73,37,17,17,25,20,20,49,63,40,19,19,15,14,19,30,52,38,17,23,15,11,18,17,41,46,19,17,16,12,14,12,21,44,23,17,19,19,17,13,15,43,23,16,17,17,13,11,11,46,26,21,17,17,17,12,10);
		wait for 10 ns;
		t_blur_matrix_int <= (92,99,107,116,116,117,112,109,84,90,102,111,118,115,115,112,70,87,96,103,115,115,115,114,60,70,97,100,110,118,116,114,43,63,85,92,103,109,115,115,30,50,69,85,96,103,111,117,17,34,57,73,86,95,105,111,11,17,34,58,70,86,118,145);
		wait for 10 ns;
		t_blur_matrix_int <= (110,108,109,107,111,113,114,112,111,109,108,107,110,112,113,114,110,107,106,113,111,109,113,116,112,108,108,107,109,113,116,116,110,107,107,105,106,116,113,117,113,107,105,108,106,113,114,117,112,106,105,104,110,112,116,119,159,162,139,104,109,132,122,119);
		wait for 10 ns;
		t_blur_matrix_int <= (115,118,121,122,116,78,26,21,116,120,122,120,94,41,16,13,117,120,123,106,56,14,10,14,122,124,115,80,20,16,14,15,121,122,100,39,16,17,17,21,122,108,61,19,19,17,17,18,119,82,25,16,17,18,17,19,98,37,16,18,16,22,17,20);
		wait for 10 ns;
		t_blur_matrix_int <= (10,11,16,16,23,27,28,34,12,13,15,22,26,34,29,29,13,16,16,19,26,28,29,31,15,18,22,22,32,27,24,23,19,19,23,24,25,30,24,26,20,17,24,27,25,27,33,27,28,24,28,21,22,30,24,27,26,25,37,24,22,28,29,26);
		wait for 10 ns;
		t_blur_matrix_int <= (27,23,27,17,18,14,17,28,28,28,24,18,15,21,20,30,28,25,26,20,16,20,30,28,29,27,18,19,24,28,30,31,34,25,21,20,27,31,21,17,28,21,21,22,27,28,25,19,25,17,25,28,30,26,24,24,26,26,23,30,29,19,24,26);
		wait for 10 ns;
		t_blur_matrix_int <= (30,26,17,21,29,29,29,32,29,19,20,20,28,28,25,30,22,18,27,19,30,30,32,30,20,20,34,24,24,27,28,27,17,22,24,28,36,25,25,26,24,27,27,21,25,20,28,37,25,29,30,26,20,19,27,60,28,32,23,20,12,18,41,84);
		wait for 10 ns;
		t_blur_matrix_int <= (42,39,33,51,72,100,114,123,34,34,40,59,91,113,122,122,32,35,58,81,110,119,120,120,31,52,84,108,122,119,118,122,39,78,107,123,122,120,120,113,62,98,121,129,124,114,110,112,95,121,128,123,120,113,109,125,115,126,124,120,111,112,121,136);
		wait for 10 ns;
		t_blur_matrix_int <= (126,126,119,116,125,135,142,145,127,129,117,124,140,148,144,145,129,122,120,137,144,147,145,145,119,119,133,143,148,147,148,140,115,127,136,148,146,148,145,144,126,138,142,146,145,147,147,144,133,141,144,143,142,143,146,146,140,139,145,142,142,142,141,140);
		wait for 10 ns;
		t_blur_matrix_int <= (60,63,58,58,59,62,60,62,58,65,58,57,57,55,53,56,55,60,57,58,57,59,56,60,67,57,59,58,57,53,55,57,54,58,55,57,60,62,59,61,57,57,58,60,59,59,59,63,62,58,60,60,57,59,58,64,61,58,62,59,61,61,63,61);
		wait for 10 ns;
		t_blur_matrix_int <= (58,58,47,53,61,78,99,112,52,51,51,49,63,78,94,110,60,57,50,52,61,77,91,110,55,53,50,51,57,73,96,104,62,59,56,50,60,80,95,106,63,55,59,52,62,78,91,105,60,57,54,51,60,77,90,106,62,63,60,53,63,75,93,104);
		wait for 10 ns;
		t_blur_matrix_int <= (120,129,135,138,139,139,139,138,120,127,133,138,142,136,138,136,118,128,137,139,141,137,140,139,119,129,136,139,137,137,138,138,117,128,134,140,141,139,138,137,118,128,136,138,142,143,142,142,118,125,137,141,143,144,142,141,116,127,136,147,143,142,145,140);
		wait for 10 ns;
		t_blur_matrix_int <= (138,138,137,125,113,98,82,69,137,137,136,121,112,99,91,75,137,137,133,120,111,99,83,66,137,140,134,121,111,100,84,67,137,137,132,124,112,95,85,66,137,135,132,125,112,98,82,59,141,138,131,124,112,99,79,64,141,141,130,123,114,98,83,68);
		wait for 10 ns;
		t_blur_matrix_int <= (52,45,43,50,54,55,61,61,55,44,44,46,49,58,60,59,57,36,39,46,48,55,53,56,46,39,40,46,50,50,55,58,46,38,38,43,48,52,57,57,50,37,39,40,44,51,60,64,44,47,43,47,42,53,57,61,48,39,42,44,47,53,59,62);
		wait for 10 ns;
		t_blur_matrix_int <= (58,61,59,65,66,69,73,66,58,62,63,64,66,63,67,65,58,58,62,59,63,65,63,62,60,60,64,65,61,64,62,60,59,67,62,63,64,65,64,66,57,62,64,65,66,68,66,62,64,66,68,65,64,66,63,65,63,68,64,63,66,69,66,67);
		wait for 10 ns;
		t_blur_matrix_int <= (68,69,69,77,75,72,76,81,62,70,72,78,72,75,73,76,68,66,68,71,68,71,72,76,64,66,67,73,70,72,72,71,66,64,65,68,72,70,70,75,64,66,64,70,70,74,68,68,64,67,63,68,69,70,74,71,67,67,68,68,69,72,75,79);
		wait for 10 ns;
		t_blur_matrix_int <= (75,80,82,81,76,76,72,80,74,80,77,76,75,75,68,95,75,78,76,78,73,65,66,147,72,76,75,77,70,66,77,187,75,78,80,74,75,63,100,205,75,79,77,77,71,65,136,205,75,79,84,87,69,71,175,199,76,78,78,80,72,79,189,188);
		wait for 10 ns;
		t_blur_matrix_int <= (170,175,97,63,73,72,70,70,196,158,89,62,70,72,69,71,200,139,80,62,71,68,67,74,183,124,81,66,63,67,71,72,169,141,88,68,65,70,70,75,169,117,75,68,64,66,68,75,159,112,70,62,66,70,70,70,158,110,64,57,62,71,68,73);
		wait for 10 ns;
		t_blur_matrix_int <= (72,77,72,80,77,79,79,79,71,78,77,80,78,77,74,71,74,75,81,84,73,78,80,77,75,77,76,80,80,80,81,83,77,70,79,83,75,81,81,87,68,73,81,88,74,79,79,85,72,76,79,86,69,76,90,74,73,79,79,64,63,87,78,87);
		wait for 10 ns;
		t_blur_matrix_int <= (82,86,89,82,91,96,94,99,78,87,84,91,92,93,102,98,81,87,84,79,97,97,99,103,85,88,89,89,93,98,102,94,83,90,81,97,96,94,103,97,84,79,96,91,102,105,88,85,84,94,98,101,97,88,96,89,91,97,93,97,91,90,79,86);
		wait for 10 ns;
		t_blur_matrix_int <= (105,104,115,103,102,105,105,104,104,103,99,109,118,112,108,105,110,106,102,101,114,106,91,101,110,103,99,108,92,93,105,108,92,104,98,78,96,108,105,107,99,80,77,100,103,108,101,99,80,91,98,104,102,95,92,98,93,106,114,94,83,96,101,85);
		wait for 10 ns;
		t_blur_matrix_int <= (109,108,108,113,112,108,98,94,100,109,108,112,95,80,95,91,107,110,107,91,84,91,88,83,110,102,91,93,87,71,72,107,97,89,103,82,76,77,110,147,97,91,81,76,80,123,141,143,81,80,75,73,131,148,156,154,80,76,85,127,139,154,159,167);
		wait for 10 ns;
		t_blur_matrix_int <= (98,80,78,96,152,167,168,170,87,80,116,145,142,171,178,180,91,122,156,160,154,173,186,176,140,145,149,172,170,160,176,155,155,157,165,175,151,144,157,162,165,165,161,155,145,138,144,155,167,157,149,143,146,145,151,165,152,142,140,143,151,163,150,146);
		wait for 10 ns;
		t_blur_matrix_int <= (175,174,182,177,166,174,168,181,164,173,163,169,179,179,185,161,168,153,156,161,176,183,170,158,161,163,161,164,162,153,164,179,157,163,171,145,148,156,175,172,179,162,147,166,164,168,154,167,144,145,166,175,172,164,156,154,165,167,158,163,166,165,163,174);
		wait for 10 ns;
		t_blur_matrix_int <= (176,171,160,163,180,189,191,183,148,152,173,178,181,183,186,189,167,178,172,178,177,186,184,186,178,174,174,166,179,185,186,183,175,170,175,179,173,184,183,180,168,179,181,173,182,179,183,173,181,178,184,175,171,176,171,183,167,187,174,184,174,170,167,173);
		wait for 10 ns;
		t_blur_matrix_int <= (190,190,184,182,190,191,196,199,186,187,193,184,188,192,187,197,192,180,187,189,186,188,187,186,184,186,178,189,184,184,187,190,187,183,187,177,187,178,183,178,181,186,185,185,177,177,170,174,172,182,186,180,165,171,190,186,183,168,162,163,178,191,190,192);
		wait for 10 ns;
		t_blur_matrix_int <= (199,194,192,197,198,195,198,197,194,194,191,196,192,194,187,189,195,196,189,187,186,188,199,198,189,185,178,187,189,193,197,200,176,181,190,197,193,194,195,197,188,193,191,192,192,193,196,196,186,190,191,188,185,187,194,193,184,185,188,189,180,175,187,195);
		wait for 10 ns;
		t_blur_matrix_int <= (193,180,192,196,198,204,206,202,197,199,192,194,199,199,200,206,195,202,200,188,194,200,200,201,196,194,201,199,192,196,199,202,197,192,189,199,197,188,195,199,190,192,192,186,192,190,189,197,188,193,193,189,189,193,192,197,193,190,193,196,195,196,196,198);
		wait for 10 ns;
		t_blur_matrix_int <= (200,200,205,206,206,208,213,220,202,194,203,204,205,209,210,221,205,199,202,204,203,205,208,210,201,201,203,201,201,204,205,207,200,199,201,198,194,197,200,202,200,197,195,201,200,200,205,200,200,201,199,203,204,202,202,201,203,199,196,198,196,195,197,198);
		wait for 10 ns;
		t_blur_matrix_int <= (223,223,176,34,31,48,70,87,223,222,209,67,28,50,65,85,221,219,219,125,29,41,63,82,214,222,223,188,50,40,57,79,211,220,222,215,128,39,51,79,204,212,221,220,199,79,45,72,201,208,212,216,217,163,53,67,200,201,203,209,215,205,101,65);
		wait for 10 ns;
		t_blur_matrix_int <= (98,107,120,121,120,120,125,124,102,109,117,121,120,122,124,124,99,108,118,122,122,125,126,125,94,106,115,120,123,123,127,122,93,108,124,123,125,124,127,129,92,106,110,131,126,126,127,129,91,105,115,129,128,127,131,128,89,104,116,124,127,126,127,127);
		wait for 10 ns;
		t_blur_matrix_int <= (122,126,125,126,110,98,88,69,123,125,120,124,111,97,89,65,126,126,123,121,113,99,85,73,122,127,124,123,113,100,81,66,126,123,125,124,115,99,82,66,126,123,123,118,111,98,84,60,129,126,128,122,108,98,77,60,126,128,125,116,111,89,71,58);
		wait for 10 ns;
		t_blur_matrix_int <= (42,27,18,15,17,16,13,16,48,23,18,17,20,17,16,10,47,23,20,18,16,14,12,12,41,23,17,16,15,10,15,17,44,20,18,14,17,15,18,77,29,13,15,12,13,30,105,194,26,14,12,16,40,137,196,209,22,14,19,61,158,207,210,185);
		wait for 10 ns;
		t_blur_matrix_int <= (12,9,18,42,84,160,192,206,11,11,26,106,189,209,216,208,19,30,124,200,213,209,192,178,52,153,203,217,200,174,182,201,171,207,213,189,155,186,207,213,208,202,169,147,195,209,213,213,196,155,155,193,211,216,210,206,143,162,199,210,213,212,207,203);
		wait for 10 ns;
		t_blur_matrix_int <= (212,209,196,160,174,196,148,109,192,186,193,205,208,212,214,143,187,201,206,212,215,218,210,196,210,216,223,223,225,228,224,221,215,221,219,217,218,223,229,229,211,212,211,210,215,216,223,231,205,206,210,205,199,208,219,230,203,204,201,198,198,209,216,227);
		wait for 10 ns;
		t_blur_matrix_int <= (56,18,19,14,21,24,21,23,26,14,18,20,19,28,18,25,43,14,21,20,21,22,22,26,104,16,21,20,23,19,26,34,171,22,21,21,21,21,22,25,203,40,21,18,17,23,25,27,212,67,21,18,19,22,21,25,219,77,19,17,18,19,22,25);
		wait for 10 ns;
		t_blur_matrix_int <= (28,24,27,28,23,32,34,31,32,23,27,25,25,29,34,27,34,28,29,38,31,23,27,26,29,24,23,31,30,29,24,25,29,27,29,22,24,21,20,23,28,28,27,24,24,22,24,28,23,27,29,24,20,25,20,19,25,28,30,19,19,21,21,18);
		wait for 10 ns;
		t_blur_matrix_int <= (27,29,24,27,20,21,26,30,25,29,30,21,20,24,25,31,27,27,30,27,20,26,35,39,25,26,26,25,27,27,26,28,23,23,21,24,28,30,25,25,25,18,26,25,26,24,28,25,15,18,28,25,30,31,27,26,14,21,22,20,27,28,27,20);
		wait for 10 ns;
		t_blur_matrix_int <= (27,22,22,21,16,33,73,110,24,19,13,22,36,66,103,122,27,17,18,18,53,95,119,126,25,16,16,35,81,116,128,125,21,19,36,68,105,126,127,123,20,29,56,98,119,127,127,119,22,37,81,115,130,126,121,119,26,63,106,129,130,122,120,120);
		wait for 10 ns;
		t_blur_matrix_int <= (125,126,118,111,111,119,131,140,126,121,117,112,120,130,138,143,125,117,117,114,129,137,145,149,118,116,115,126,135,143,145,146,116,117,123,134,138,141,142,141,113,121,132,139,139,141,137,141,119,129,138,137,139,139,135,138,125,135,138,138,134,136,135,137);
		wait for 10 ns;
		t_blur_matrix_int <= (139,142,140,139,136,138,138,141,144,142,138,140,138,140,137,139,139,140,141,139,137,136,138,136,139,142,136,139,138,135,139,137,138,141,140,140,139,140,135,136,140,140,137,137,138,136,138,137,139,140,139,139,136,139,138,134,138,136,137,134,137,137,136,138);
		wait for 10 ns;
		t_blur_matrix_int <= (60,61,62,64,60,65,66,63,60,63,63,62,65,64,68,64,63,68,65,62,64,68,64,63,66,65,65,68,65,65,69,68,70,67,66,67,69,63,66,67,66,67,69,69,67,67,66,65,67,69,65,62,64,63,67,67,69,66,66,64,63,63,66,66);
		wait for 10 ns;
		t_blur_matrix_int <= (65,62,65,61,63,80,93,102,64,62,63,60,63,78,89,109,62,60,62,56,66,74,95,105,65,63,59,63,63,72,93,105,66,62,64,59,66,79,91,107,68,64,63,65,70,79,92,108,69,58,66,63,73,77,95,108,70,63,61,64,70,78,95,108);
		wait for 10 ns;
		t_blur_matrix_int <= (117,130,136,141,146,143,146,143,116,126,138,141,145,143,146,143,117,129,135,142,140,143,142,146,120,128,134,141,142,142,144,140,119,128,134,138,143,143,148,146,119,123,130,142,140,145,149,148,120,127,134,141,144,147,147,149,123,132,139,139,147,151,150,148);
		wait for 10 ns;
		t_blur_matrix_int <= (143,140,135,127,116,101,82,69,140,143,134,129,119,101,82,69,144,144,139,126,118,103,82,67,143,146,137,129,117,105,86,66,143,142,140,131,120,105,85,73,146,147,147,128,120,103,87,69,147,147,145,134,122,105,88,69,150,150,147,136,122,105,87,66);
		wait for 10 ns;
		t_blur_matrix_int <= (52,42,46,45,49,55,58,61,52,46,43,47,52,56,61,62,50,43,44,46,53,60,64,63,50,42,47,48,52,52,61,60,50,41,44,47,54,52,59,64,47,46,44,47,54,59,60,61,52,42,41,48,56,62,58,64,49,47,45,51,58,59,59,60);
		wait for 10 ns;
		t_blur_matrix_int <= (62,62,63,67,66,70,65,63,65,67,65,68,67,63,67,67,67,67,61,72,69,66,67,74,64,65,65,66,65,67,72,70,69,70,68,67,67,69,62,71,63,63,65,68,69,68,63,69,66,69,64,68,67,64,68,68,69,64,63,69,66,67,66,64);
		wait for 10 ns;
		t_blur_matrix_int <= (63,68,72,71,72,72,74,74,66,64,69,73,69,70,76,76,69,64,68,72,75,76,75,74,67,65,64,68,79,74,75,78,66,62,65,65,72,71,72,78,68,65,63,67,67,71,74,73,67,66,65,69,67,73,71,74,59,65,67,70,69,74,72,75);
		wait for 10 ns;
		t_blur_matrix_int <= (77,78,81,70,63,90,206,185,77,79,77,72,66,112,205,186,82,79,79,70,62,146,201,189,76,79,80,69,66,169,202,177,76,79,73,64,64,192,200,158,77,74,71,60,76,204,188,137,71,74,70,60,97,209,190,131,71,70,65,54,130,209,179,143);
		wait for 10 ns;
		t_blur_matrix_int <= (149,123,72,58,71,68,72,76,146,95,75,63,71,62,73,71,122,92,73,60,61,64,67,66,112,82,78,64,62,62,68,71,102,84,81,69,59,67,70,72,103,98,87,70,73,65,69,74,114,93,88,71,69,71,74,65,113,94,93,66,72,71,70,75);
		wait for 10 ns;
		t_blur_matrix_int <= (71,72,62,71,79,84,88,88,68,56,73,84,85,79,89,96,63,75,79,86,76,90,78,84,75,77,72,75,80,64,75,93,74,71,67,75,65,75,85,84,61,72,64,59,78,79,85,84,68,62,62,78,63,78,73,64,75,72,69,66,77,79,74,82);
		wait for 10 ns;
		t_blur_matrix_int <= (92,93,83,94,89,78,90,95,84,91,91,82,95,94,82,91,97,82,71,90,86,89,94,96,78,73,93,92,88,94,93,95,86,87,83,88,91,98,97,88,72,79,94,93,96,88,75,84,82,88,83,89,82,73,87,92,82,90,89,79,81,94,93,90);
		wait for 10 ns;
		t_blur_matrix_int <= (95,103,100,93,98,105,95,81,104,99,113,110,103,95,74,67,103,99,91,93,95,72,60,99,90,82,88,95,76,71,101,123,85,93,87,78,77,105,122,141,90,84,82,76,107,111,128,132,83,82,86,114,121,119,123,126,84,79,115,128,118,128,114,114);
		wait for 10 ns;
		t_blur_matrix_int <= (71,89,138,139,139,158,155,148,96,119,133,154,146,140,136,138,137,139,128,139,156,125,119,129,130,140,142,117,121,132,120,141,133,134,131,117,112,115,154,120,137,116,119,119,132,128,103,120,124,116,117,129,136,100,121,137,113,116,141,110,98,119,129,134);
		wait for 10 ns;
		t_blur_matrix_int <= (147,137,132,154,163,139,151,164,137,151,158,135,134,150,170,165,154,161,131,136,152,156,154,171,145,123,140,160,158,150,151,154,108,141,152,155,155,155,161,165,135,137,149,151,154,162,161,159,145,142,127,152,166,160,157,145,135,141,148,145,153,156,151,150);
		wait for 10 ns;
		t_blur_matrix_int <= (166,169,161,156,158,171,177,176,165,161,164,157,170,171,179,167,160,157,173,172,160,158,165,175,167,171,163,178,160,156,159,163,157,162,159,153,165,161,154,168,151,146,148,154,152,177,173,157,147,147,145,143,169,166,175,166,145,146,159,161,141,169,154,145);
		wait for 10 ns;
		t_blur_matrix_int <= (170,165,177,169,180,174,179,165,172,171,163,175,167,178,162,151,167,165,168,161,176,151,148,154,171,164,167,167,146,143,162,170,161,174,164,143,139,157,178,174,164,148,144,153,168,163,158,172,138,130,154,171,160,157,162,154,128,149,165,161,156,159,155,163);
		wait for 10 ns;
		t_blur_matrix_int <= (160,157,173,183,179,184,188,189,153,162,185,172,177,180,187,189,166,178,181,175,166,172,181,182,165,164,179,176,176,167,178,180,169,163,171,179,179,172,171,181,173,165,168,161,159,177,174,158,172,171,160,162,163,154,165,171,158,161,167,152,172,163,151,169);
		wait for 10 ns;
		t_blur_matrix_int <= (191,181,182,191,190,186,178,189,188,187,180,179,188,189,187,182,186,188,187,186,186,184,189,190,180,185,186,178,189,195,187,188,178,175,183,175,184,191,193,191,167,179,181,181,181,191,195,192,157,166,183,186,180,170,176,166,174,171,179,158,151,142,159,162);
		wait for 10 ns;
		t_blur_matrix_int <= (194,193,189,191,194,201,196,190,190,195,192,187,179,186,167,182,183,194,198,185,148,148,179,193,192,191,183,157,147,169,183,186,192,185,142,147,177,184,181,184,171,154,164,172,178,178,185,188,152,172,178,183,177,177,172,175,172,180,169,165,163,172,173,178);
		wait for 10 ns;
		t_blur_matrix_int <= (191,185,189,197,197,199,196,200,190,185,193,196,196,197,192,200,193,190,191,197,192,195,193,193,191,192,194,197,192,194,195,194,189,193,190,193,193,194,193,192,190,188,188,187,184,190,188,189,183,180,186,189,186,182,184,181,186,180,185,190,187,178,173,181);
		wait for 10 ns;
		t_blur_matrix_int <= (199,202,201,204,210,214,182,103,198,198,200,199,205,208,210,191,195,197,194,194,199,207,207,211,191,189,188,192,195,198,204,207,192,191,189,185,190,192,195,200,190,190,190,189,182,188,188,189,180,187,189,188,181,179,186,180,179,179,184,182,181,172,178,177);
		wait for 10 ns;
		t_blur_matrix_int <= (87,98,116,121,125,126,129,127,136,98,111,122,122,125,128,126,206,141,106,118,121,123,123,125,209,194,125,118,127,126,123,120,200,205,161,116,127,124,121,116,200,201,191,120,122,125,120,117,186,194,195,131,121,122,120,119,180,185,192,167,113,119,133,176);
		wait for 10 ns;
		t_blur_matrix_int <= (127,126,120,115,103,81,65,45,126,124,120,116,97,79,53,38,123,121,118,109,91,73,69,121,120,120,111,101,94,115,172,207,121,116,109,126,172,201,208,192,112,119,158,195,208,198,178,181,143,177,201,205,182,178,181,169,193,200,184,182,188,179,177,193);
		wait for 10 ns;
		t_blur_matrix_int <= (21,35,102,182,210,204,179,150,73,155,201,210,190,169,163,192,188,211,196,182,167,171,193,208,212,189,179,178,181,200,208,205,177,179,170,188,201,206,205,203,180,173,194,202,206,203,200,198,183,201,205,201,199,196,192,193,203,205,198,198,195,191,192,194);
		wait for 10 ns;
		t_blur_matrix_int <= (175,200,210,208,207,206,205,197,205,211,207,204,203,201,198,193,207,206,201,201,200,197,195,191,206,201,196,197,197,191,192,193,201,195,194,197,191,192,194,195,196,193,195,190,196,196,195,196,192,192,193,196,196,198,194,198,194,193,194,196,197,195,197,196);
		wait for 10 ns;
		t_blur_matrix_int <= (187,196,196,199,205,211,216,226,194,195,195,202,207,213,219,222,193,196,199,207,210,213,218,221,197,199,200,206,211,214,216,219,196,201,206,209,210,214,216,220,202,205,208,208,212,216,216,218,199,204,206,207,213,216,217,219,195,200,203,208,214,215,217,218);
		wait for 10 ns;
		t_blur_matrix_int <= (221,75,17,16,22,23,31,30,218,67,14,17,21,25,30,35,212,57,22,23,24,26,24,28,205,35,24,14,19,21,20,24,184,20,20,26,27,26,22,22,152,20,18,21,27,23,24,22,117,20,25,33,30,28,26,25,81,27,24,26,26,30,28,25);
		wait for 10 ns;
		t_blur_matrix_int <= (27,19,17,15,17,24,18,19,31,20,23,17,16,17,15,20,32,21,25,20,20,22,15,26,33,33,31,21,19,17,23,27,23,26,24,17,14,19,17,25,25,25,24,20,19,18,15,24,24,22,19,18,13,18,19,26,24,22,17,12,18,27,20,26);
		wait for 10 ns;
		t_blur_matrix_int <= (21,20,22,27,25,20,17,22,22,26,23,22,19,12,10,30,28,26,31,26,12,6,15,52,22,26,25,19,7,10,31,82,23,25,26,18,9,20,56,103,25,21,22,18,20,46,89,121,25,30,26,31,35,72,109,123,24,32,33,39,55,92,121,124);
		wait for 10 ns;
		t_blur_matrix_int <= (42,91,124,132,127,122,116,126,68,116,131,126,120,119,121,133,102,123,129,124,118,119,127,138,116,132,130,123,116,128,134,139,127,131,124,121,124,131,139,142,129,128,122,119,125,135,140,140,128,122,121,121,133,137,137,141,120,118,119,128,135,141,136,136);
		wait for 10 ns;
		t_blur_matrix_int <= (136,138,138,137,139,135,137,136,139,143,140,138,137,135,137,136,137,139,140,135,136,136,134,136,138,140,137,136,136,135,134,133,136,141,141,135,136,135,136,133,139,136,138,136,136,136,133,137,139,139,133,136,134,139,136,137,138,138,140,135,135,134,135,136);
		wait for 10 ns;
		t_blur_matrix_int <= (139,134,139,133,135,133,138,137,138,139,134,135,132,129,136,134,135,133,136,138,134,134,135,134,137,134,133,134,132,132,131,134,139,135,131,135,130,131,133,130,135,135,136,134,133,131,132,132,134,132,134,132,134,131,133,128,136,134,133,131,132,131,132,131);
		wait for 10 ns;
		t_blur_matrix_int <= (66,70,65,64,67,67,67,64,64,65,67,68,68,65,60,66,70,64,66,65,68,57,64,65,70,65,62,67,67,64,62,64,66,60,65,67,68,66,64,65,60,67,70,62,61,63,63,64,64,63,64,67,62,63,62,63,64,65,62,68,59,64,65,64);
		wait for 10 ns;
		t_blur_matrix_int <= (69,64,64,61,66,80,93,108,68,63,63,65,72,81,96,108,68,64,67,65,72,82,93,107,62,62,63,63,69,80,92,110,64,64,63,60,67,77,92,109,64,69,63,63,67,82,92,110,61,64,61,63,71,77,96,110,63,62,62,65,66,78,98,110);
		wait for 10 ns;
		t_blur_matrix_int <= (121,133,138,143,146,145,149,151,123,128,140,143,149,149,153,153,120,133,141,146,149,149,155,151,119,129,142,148,150,153,154,150,118,133,140,144,153,149,152,148,119,133,141,146,151,149,153,150,122,133,141,150,151,150,151,152,126,134,144,149,147,147,152,149);
		wait for 10 ns;
		t_blur_matrix_int <= (149,151,146,139,122,109,84,70,151,149,146,135,122,108,86,72,151,151,145,136,123,106,81,73,150,152,144,135,120,104,83,74,151,150,146,138,118,106,92,72,148,153,145,134,122,108,88,74,147,149,145,134,124,105,88,70,145,149,141,136,121,107,91,71);
		wait for 10 ns;
		t_blur_matrix_int <= (53,43,46,50,62,63,56,60,51,44,41,45,53,55,58,63,52,43,42,47,52,54,62,58,51,39,41,45,54,56,62,64,51,44,43,46,51,58,61,63,55,44,46,52,59,57,62,58,50,46,42,51,56,62,62,62,54,48,45,46,54,62,63,62);
		wait for 10 ns;
		t_blur_matrix_int <= (63,69,68,66,64,65,64,65,57,64,65,70,63,65,62,63,60,61,64,71,66,63,62,66,62,64,61,65,64,62,64,65,60,65,62,65,63,66,65,64,61,66,66,68,64,61,66,67,63,63,72,67,66,63,62,66,69,67,63,63,66,63,65,64);
		wait for 10 ns;
		t_blur_matrix_int <= (60,64,70,65,68,69,69,70,62,67,63,64,66,68,69,74,65,63,67,64,63,69,72,68,63,62,63,66,67,69,73,70,63,67,63,63,69,67,67,72,60,67,62,63,69,68,70,72,63,64,61,67,66,67,65,68,64,64,64,68,66,66,71,64);
		wait for 10 ns;
		t_blur_matrix_int <= (71,67,59,57,156,205,181,143,70,65,57,60,188,205,171,152,66,65,55,70,205,199,175,158,65,70,54,76,207,196,167,161,67,65,56,84,212,191,172,154,67,65,53,92,213,194,168,150,66,64,54,86,211,180,166,152,66,63,55,95,213,181,173,144);
		wait for 10 ns;
		t_blur_matrix_int <= (125,104,92,80,64,69,67,74,119,105,91,75,72,68,78,75,121,120,91,92,76,85,75,66,124,112,105,96,92,85,78,82,115,121,103,106,81,106,84,77,148,126,112,113,96,93,90,70,136,137,118,112,110,106,89,82,137,128,124,112,111,99,103,92);
		wait for 10 ns;
		t_blur_matrix_int <= (73,71,68,81,64,80,76,73,70,65,74,72,78,80,83,83,69,68,73,75,74,80,81,79,71,72,71,70,78,75,63,81,66,71,66,78,70,71,74,82,72,73,67,69,72,81,71,91,79,73,49,65,74,68,84,87,78,64,66,60,58,77,82,78);
		wait for 10 ns;
		t_blur_matrix_int <= (89,86,75,84,89,96,93,79,82,78,83,88,95,88,77,74,87,97,86,92,96,79,71,104,83,83,93,89,85,79,95,112,88,84,79,79,77,98,114,105,92,70,65,71,107,119,104,114,82,71,69,98,115,115,108,102,77,70,106,107,110,110,109,100);
		wait for 10 ns;
		t_blur_matrix_int <= (75,106,119,121,124,130,113,103,107,123,114,123,126,117,111,113,116,124,121,114,109,112,120,124,117,123,120,107,104,117,138,94,119,121,108,110,116,128,89,89,117,107,114,113,127,84,91,109,109,109,127,113,80,86,115,118,106,119,121,81,86,106,112,121);
		wait for 10 ns;
		t_blur_matrix_int <= (116,133,112,97,116,125,138,132,119,110,98,112,124,124,120,141,96,95,112,120,119,125,126,128,103,117,127,121,121,126,137,115,112,123,124,122,129,134,121,102,120,117,121,128,130,127,111,107,123,122,121,130,118,124,114,124,120,128,120,114,114,115,131,132);
		wait for 10 ns;
		t_blur_matrix_int <= (129,147,153,131,129,141,148,151,149,138,132,144,136,139,140,162,147,124,126,133,141,145,156,145,111,133,121,139,156,157,153,156,112,111,135,141,143,166,152,147,120,125,121,138,134,134,157,130,133,138,113,111,146,131,117,125,114,119,121,115,125,125,118,137);
		wait for 10 ns;
		t_blur_matrix_int <= (159,152,150,166,154,131,136,136,166,168,148,144,148,128,151,162,157,164,157,130,128,142,155,169,141,133,135,132,159,161,142,152,137,111,138,163,159,159,154,140,124,138,152,153,161,156,148,147,145,158,157,146,143,143,154,149,148,151,154,149,143,141,140,152);
		wait for 10 ns;
		t_blur_matrix_int <= (164,160,154,160,163,162,163,153,156,161,156,149,155,168,160,155,160,145,156,158,150,150,164,155,154,149,153,156,167,154,144,162,140,160,155,154,161,168,153,148,142,143,159,158,156,156,162,151,147,146,138,150,159,150,140,141,148,153,148,134,143,155,144,139);
		wait for 10 ns;
		t_blur_matrix_int <= (158,158,153,167,157,168,167,168,161,154,150,157,168,156,176,185,159,155,152,147,152,168,166,167,158,155,159,149,156,148,161,159,160,157,154,152,142,153,150,155,140,130,148,164,149,140,149,161,147,142,142,139,151,156,152,142,147,144,149,149,141,144,130,132);
		wait for 10 ns;
		t_blur_matrix_int <= (179,175,178,154,153,170,174,172,177,167,161,165,167,163,166,170,164,165,168,169,169,170,171,164,159,173,177,170,163,166,168,157,167,166,165,162,158,168,171,169,156,161,144,154,164,162,171,174,141,147,160,153,157,163,159,174,144,150,157,158,156,158,154,156);
		wait for 10 ns;
		t_blur_matrix_int <= (179,172,159,164,180,180,186,178,180,181,179,172,175,183,184,181,165,175,178,184,175,177,181,179,166,174,173,183,180,172,176,177,159,167,174,181,181,179,166,161,173,157,171,178,174,171,165,158,173,170,161,167,168,160,161,157,174,171,165,158,159,162,158,156);
		wait for 10 ns;
		t_blur_matrix_int <= (188,184,180,185,181,172,170,176,178,182,177,164,176,169,169,173,177,169,169,169,155,163,171,174,169,169,161,156,160,156,167,174,165,168,173,163,154,162,151,170,160,165,163,172,166,152,162,151,150,166,168,168,165,150,153,137,150,148,163,171,158,153,133,136);
		wait for 10 ns;
		t_blur_matrix_int <= (179,178,174,180,177,173,175,182,176,176,170,176,174,172,162,175,175,164,174,169,172,164,154,155,173,170,160,160,163,149,143,153,169,168,151,159,137,146,162,190,165,159,144,143,149,187,196,185,155,145,148,168,194,192,167,171,138,162,186,189,167,169,178,180);
		wait for 10 ns;
		t_blur_matrix_int <= (175,176,182,190,143,154,190,206,171,175,175,184,185,196,198,184,170,169,182,193,191,176,173,189,175,196,194,171,165,166,186,188,194,179,157,164,186,185,190,196,171,169,182,177,186,193,198,197,183,180,185,193,197,194,194,192,185,191,197,199,191,189,189,187);
		wait for 10 ns;
		t_blur_matrix_int <= (193,170,178,177,179,192,198,200,182,184,183,187,194,201,197,196,185,184,194,201,204,199,194,188,188,196,202,205,200,195,184,187,198,199,198,198,193,187,188,191,195,192,193,192,188,188,189,192,188,183,185,185,188,190,187,192,181,181,180,184,188,186,192,190);
		wait for 10 ns;
		t_blur_matrix_int <= (200,197,196,195,192,193,191,193,196,196,193,193,191,191,188,192,191,194,193,192,191,191,189,194,193,190,193,192,186,189,191,194,191,194,191,191,191,191,195,195,192,190,190,191,190,193,196,196,191,192,187,195,195,192,195,197,193,192,190,193,191,197,195,199);
		wait for 10 ns;
		t_blur_matrix_int <= (192,194,198,199,197,195,193,191,192,196,196,197,194,196,187,186,195,198,195,196,197,186,177,184,193,197,196,198,191,168,159,177,197,195,198,198,165,149,149,165,195,197,197,176,148,137,140,155,200,192,191,155,138,136,139,164,198,199,163,138,132,146,164,163);
		wait for 10 ns;
		t_blur_matrix_int <= (193,202,205,207,214,216,219,214,195,203,202,204,215,218,220,196,195,201,202,206,214,216,216,155,190,198,199,202,209,212,213,94,181,198,195,198,209,209,201,44,183,181,176,187,202,207,148,16,163,128,158,183,195,206,76,18,106,122,158,179,194,181,23,21);
		wait for 10 ns;
		t_blur_matrix_int <= (54,17,26,26,24,31,23,28,27,17,19,17,21,17,23,35,15,11,17,20,22,17,24,23,16,11,18,20,19,27,20,30,16,15,16,17,17,25,23,36,17,20,20,19,24,24,18,25,17,33,30,25,21,30,26,24,12,27,34,32,28,25,18,17);
		wait for 10 ns;
		t_blur_matrix_int <= (29,20,22,17,21,23,18,24,30,24,17,14,23,23,20,29,19,16,16,22,22,26,30,27,29,20,20,16,21,31,27,19,37,16,23,21,28,31,28,16,22,18,21,19,21,22,27,24,20,14,21,19,13,23,39,47,19,19,26,16,22,32,45,57);
		wait for 10 ns;
		t_blur_matrix_int <= (27,28,36,48,80,114,123,124,35,37,48,72,102,122,125,119,21,36,58,92,115,127,125,119,17,41,77,110,125,125,120,117,19,50,98,124,131,121,118,121,33,73,111,127,126,120,118,127,57,100,121,128,120,119,120,130,88,115,124,124,118,118,127,136);
		wait for 10 ns;
		t_blur_matrix_int <= (121,118,124,132,138,140,139,136,118,121,131,137,140,139,141,138,118,125,134,137,142,140,139,138,122,128,137,138,140,140,139,138,131,138,140,137,141,140,136,139,136,140,140,142,143,141,138,135,135,139,138,139,140,136,138,138,139,139,140,140,137,132,138,138);
		wait for 10 ns;
		t_blur_matrix_int <= (138,137,136,135,135,133,137,135,138,138,137,134,135,136,134,137,138,135,135,135,135,133,136,134,137,140,140,134,135,139,136,136,141,139,137,138,134,135,137,139,138,140,139,133,136,134,137,136,135,142,137,134,140,135,140,135,138,137,136,139,136,137,135,136);
		wait for 10 ns;
		t_blur_matrix_int <= (131,133,133,133,134,130,133,132,134,133,134,134,132,133,136,134,136,134,134,132,134,133,135,134,135,136,138,134,134,135,139,132,136,136,135,137,133,138,139,135,137,134,135,139,137,136,134,133,137,136,140,139,134,134,137,133,138,137,137,140,135,133,136,135);
		wait for 10 ns;
		t_blur_matrix_int <= (64,64,59,62,61,58,59,63,59,74,62,63,62,66,64,61,62,63,62,61,60,62,62,60,65,66,66,60,56,61,61,64,61,62,64,66,65,60,63,63,62,63,63,66,65,65,62,62,67,62,67,64,60,65,67,66,66,68,62,67,61,65,65,65);
		wait for 10 ns;
		t_blur_matrix_int <= (61,63,64,64,66,81,97,113,61,62,63,64,68,83,96,110,59,60,60,62,69,79,100,109,60,62,60,64,74,85,97,109,64,62,64,64,71,83,98,112,64,66,68,70,72,84,95,108,64,63,72,70,71,83,98,111,65,66,67,68,72,82,100,112);
		wait for 10 ns;
		t_blur_matrix_int <= (123,133,142,146,147,147,148,148,123,135,142,144,151,150,149,150,125,134,143,149,150,149,147,148,123,133,141,146,148,150,146,148,121,133,141,146,149,149,152,153,121,136,139,148,151,149,149,150,121,134,142,151,148,150,151,149,123,132,143,148,148,152,151,150);
		wait for 10 ns;
		t_blur_matrix_int <= (146,148,144,135,121,107,87,71,150,149,145,136,124,114,89,70,148,148,148,136,121,108,92,71,152,145,146,136,122,112,91,74,151,151,145,135,123,114,93,78,147,149,144,137,124,113,97,67,148,152,145,140,125,111,90,67,152,151,145,140,130,111,93,72);
		wait for 10 ns;
		t_blur_matrix_int <= (55,41,46,46,52,61,58,64,54,41,44,48,56,61,61,65,59,44,48,48,54,58,62,65,50,43,45,50,57,57,60,64,58,41,47,43,53,57,61,62,53,41,39,46,52,60,62,66,53,39,39,49,52,55,59,67,54,42,36,42,57,56,61,65);
		wait for 10 ns;
		t_blur_matrix_int <= (63,68,66,64,63,65,63,65,65,67,65,65,66,59,61,65,64,62,64,63,63,60,66,62,64,66,63,63,65,63,65,63,60,66,60,62,62,57,63,64,60,66,65,62,62,60,66,65,66,61,64,59,59,60,65,62,64,62,65,64,68,62,62,68);
		wait for 10 ns;
		t_blur_matrix_int <= (64,62,64,65,69,64,68,66,64,65,64,66,69,63,65,64,63,66,69,68,66,62,68,65,59,62,62,65,64,60,66,66,65,65,65,63,62,66,65,61,62,62,66,65,64,63,64,59,63,65,59,61,67,62,65,60,63,62,59,66,64,62,58,62);
		wait for 10 ns;
		t_blur_matrix_int <= (63,62,51,107,205,175,166,150,63,56,48,123,206,175,160,154,60,55,49,146,196,170,169,153,58,54,47,157,190,182,164,175,58,50,48,175,196,184,185,155,58,46,45,171,197,189,172,189,55,47,43,171,205,185,193,161,60,47,43,169,201,197,170,194);
		wait for 10 ns;
		t_blur_matrix_int <= (141,134,144,110,105,111,108,87,137,131,113,124,108,101,112,91,156,116,137,118,107,96,112,94,144,144,118,136,116,111,106,106,169,141,146,130,126,99,120,111,148,155,138,140,113,125,109,126,170,137,152,129,141,131,123,122,153,152,135,142,125,117,132,122);
		wait for 10 ns;
		t_blur_matrix_int <= (71,68,63,56,72,75,72,68,74,71,67,73,75,74,68,69,80,82,76,67,71,65,73,105,84,89,76,74,63,67,101,95,101,75,72,59,61,102,109,104,103,97,66,52,82,98,106,104,122,90,68,71,93,95,93,96,123,94,80,90,85,91,93,94);
		wait for 10 ns;
		t_blur_matrix_int <= (64,109,116,108,104,104,100,107,100,114,110,108,104,89,105,116,116,112,110,103,101,101,107,101,107,106,103,103,105,115,88,83,87,106,100,100,115,95,87,89,101,90,105,111,92,85,98,90,98,96,112,97,78,92,91,111,94,109,92,78,87,92,106,110);
		wait for 10 ns;
		t_blur_matrix_int <= (110,114,79,91,105,108,108,120,97,90,87,96,114,119,112,114,79,96,99,116,114,112,126,107,85,94,116,116,115,117,119,110,93,116,108,108,117,121,105,116,117,113,106,107,112,107,108,102,116,114,107,111,108,114,101,86,106,112,104,100,115,89,87,103);
		wait for 10 ns;
		t_blur_matrix_int <= (127,116,115,107,115,129,117,126,117,112,110,118,114,112,103,124,105,112,120,104,105,113,125,120,108,119,94,98,107,121,126,127,104,91,93,104,122,128,114,123,91,105,103,106,129,124,113,95,99,106,115,109,107,119,91,122,97,107,113,125,99,95,116,122);
		wait for 10 ns;
		t_blur_matrix_int <= (119,137,133,123,105,125,149,130,131,130,128,110,123,122,138,145,124,112,104,125,137,143,126,131,113,102,124,129,136,131,137,122,100,122,135,135,128,129,132,124,106,121,130,140,135,122,114,93,121,117,123,119,100,68,79,92,127,126,113,83,67,91,125,110);
		wait for 10 ns;
		t_blur_matrix_int <= (136,143,136,138,152,150,140,146,135,123,129,133,140,164,144,134,134,134,128,132,139,137,140,130,119,139,145,125,125,129,116,115,125,119,139,138,139,132,126,118,100,106,104,114,119,129,123,97,87,72,69,64,78,102,108,80,105,88,90,80,75,53,62,79);
		wait for 10 ns;
		t_blur_matrix_int <= (149,146,147,138,134,130,159,148,138,134,138,145,142,142,134,151,134,135,141,138,146,151,141,129,131,136,143,146,144,135,128,125,105,98,102,84,94,134,137,138,121,121,118,85,43,126,142,135,124,120,132,120,77,94,121,126,130,145,143,140,118,95,84,82);
		wait for 10 ns;
		t_blur_matrix_int <= (140,144,151,140,125,139,148,147,150,119,125,138,154,140,139,148,121,118,144,156,142,146,147,152,142,142,137,145,145,136,140,147,142,143,140,143,136,145,136,134,138,139,134,133,132,138,138,144,139,138,141,141,115,118,122,121,90,87,95,135,136,134,141,121);
		wait for 10 ns;
		t_blur_matrix_int <= (152,150,148,159,157,150,151,147,140,148,153,148,155,149,140,154,143,136,151,148,156,147,147,140,146,142,137,148,137,146,142,148,143,149,141,132,148,137,145,144,136,142,144,132,133,136,131,139,125,141,136,140,120,106,91,55,85,112,106,120,139,93,112,53);
		wait for 10 ns;
		t_blur_matrix_int <= (160,171,163,157,147,153,157,158,148,151,155,151,155,147,152,156,149,139,136,144,156,150,139,148,134,141,142,139,141,146,136,139,144,132,145,147,123,139,132,127,139,139,131,140,129,120,131,137,130,134,134,119,128,114,150,180,31,108,135,118,119,163,179,166);
		wait for 10 ns;
		t_blur_matrix_int <= (144,154,149,162,155,142,130,147,144,147,140,144,143,144,168,188,146,126,138,129,148,180,181,164,140,127,140,173,183,174,158,161,133,164,179,181,152,158,177,171,172,191,159,157,158,173,185,183,176,158,151,169,182,185,188,191,143,151,166,182,198,194,191,182);
		wait for 10 ns;
		t_blur_matrix_int <= (176,192,169,166,171,170,177,191,176,153,159,173,175,190,192,200,160,169,173,185,192,196,193,189,168,182,192,187,187,184,183,177,184,195,194,187,180,177,172,173,186,192,189,179,178,179,182,178,186,188,181,177,180,183,183,183,182,186,185,185,182,184,182,184);
		wait for 10 ns;
		t_blur_matrix_int <= (200,195,195,193,191,185,174,183,197,194,191,185,183,184,184,185,189,185,183,184,178,185,184,185,171,171,183,179,183,186,188,188,175,176,181,184,186,185,186,189,180,184,185,187,186,188,190,190,184,185,187,190,188,192,191,189,186,187,189,193,191,191,193,192);
		wait for 10 ns;
		t_blur_matrix_int <= (185,181,181,186,187,190,193,192,183,183,186,187,189,191,193,193,187,186,188,191,191,195,193,193,187,187,193,193,196,195,196,194,190,193,194,196,195,196,195,194,192,193,194,195,195,193,196,196,194,193,193,198,195,196,196,195,192,196,196,196,194,196,196,196);
		wait for 10 ns;
		t_blur_matrix_int <= (192,193,192,196,192,201,199,199,191,194,195,195,196,198,200,202,194,196,194,196,199,201,201,202,193,195,196,198,201,202,205,197,194,196,196,201,202,203,208,170,195,198,199,203,202,205,197,135,195,199,201,204,206,202,160,144,195,200,202,206,208,174,149,134);
		wait for 10 ns;
		t_blur_matrix_int <= (200,188,134,136,142,162,166,107,200,152,134,145,161,160,113,119,182,133,133,157,157,119,126,144,141,132,150,152,117,135,151,136,130,149,145,121,140,136,101,85,148,139,130,122,84,77,62,88,136,131,89,59,49,63,72,118,104,59,52,59,59,76,96,154);
		wait for 10 ns;
		t_blur_matrix_int <= (109,137,160,180,208,118,12,13,134,154,159,181,210,65,12,16,150,137,163,203,184,23,19,19,116,127,179,217,115,20,14,18,108,157,203,210,47,13,17,21,122,181,216,172,19,14,11,20,161,208,218,94,10,10,9,19,197,213,186,26,12,12,12,20);
		wait for 10 ns;
		t_blur_matrix_int <= (13,15,24,41,36,23,15,15,14,17,24,22,26,20,16,19,21,22,23,26,22,37,16,17,23,25,24,22,26,20,34,26,23,31,27,27,33,24,33,44,27,27,24,22,24,22,28,41,22,23,22,18,19,20,27,28,25,22,23,21,18,26,24,30);
		wait for 10 ns;
		t_blur_matrix_int <= (21,25,23,17,22,35,49,73,26,23,22,18,29,46,55,94,23,24,24,21,34,43,78,110,29,27,20,31,44,55,99,124,29,22,29,20,39,73,113,127,25,29,29,32,48,96,125,128,23,26,26,37,75,110,126,127,26,27,31,50,95,121,126,124);
		wait for 10 ns;
		t_blur_matrix_int <= (109,122,127,122,119,121,132,136,123,131,122,117,118,127,137,138,130,127,119,121,121,129,135,137,128,126,116,117,127,137,136,139,126,121,118,124,131,135,137,136,121,120,122,128,135,139,139,137,118,118,126,131,137,139,137,138,120,119,130,139,139,137,137,137);
		wait for 10 ns;
		t_blur_matrix_int <= (140,141,140,143,141,134,140,134,139,143,137,137,142,137,134,136,141,138,140,137,136,134,135,132,140,140,134,137,134,131,135,137,137,136,136,134,136,135,136,132,137,137,136,136,133,133,132,133,137,136,137,134,133,136,135,133,136,140,135,135,135,134,136,135);
		wait for 10 ns;
		t_blur_matrix_int <= (136,138,138,139,140,133,134,135,137,138,137,138,138,137,136,136,134,135,139,137,135,136,137,135,136,138,136,136,134,139,135,134,133,135,138,136,135,134,136,135,136,134,133,135,133,136,135,133,133,136,134,133,134,135,132,135,134,136,134,135,131,135,134,136);
		wait for 10 ns;
		t_blur_matrix_int <= (134,136,140,138,138,134,137,134,136,133,138,136,134,135,139,137,140,136,136,133,136,134,134,135,138,137,135,135,135,135,136,136,136,138,136,135,138,135,134,133,136,136,135,136,133,134,134,133,133,139,135,137,130,133,132,133,135,133,134,133,133,129,136,130);
		wait for 10 ns;
		t_blur_matrix_int <= (67,66,61,67,68,63,63,66,63,69,66,65,61,74,64,67,66,65,69,69,69,65,68,64,63,68,69,71,70,64,67,66,67,67,69,71,68,66,65,60,66,69,68,70,70,68,63,61,73,72,71,69,72,64,61,64,71,73,75,68,70,60,66,65);
		wait for 10 ns;
		t_blur_matrix_int <= (66,63,63,66,73,84,100,111,69,70,70,71,79,90,101,113,65,70,69,70,74,83,104,114,68,63,72,72,74,85,102,113,65,75,72,69,75,86,99,113,64,70,66,70,77,88,101,112,62,67,70,71,74,85,100,114,66,65,65,68,72,89,96,113);
		wait for 10 ns;
		t_blur_matrix_int <= (123,133,143,149,150,150,157,150,125,133,143,149,154,149,152,150,126,133,145,152,150,151,153,150,125,138,147,147,154,149,149,152,125,137,149,151,146,148,151,151,125,134,146,150,153,149,149,153,122,134,143,148,148,148,150,154,122,134,142,149,152,149,150,148);
		wait for 10 ns;
		t_blur_matrix_int <= (150,151,146,138,128,112,92,72,151,152,147,137,127,111,93,72,151,152,145,140,126,111,92,76,148,153,147,136,129,114,92,74,150,151,149,139,128,111,95,70,149,149,144,140,130,111,94,70,149,149,147,139,130,112,96,69,151,149,146,139,129,114,93,72);
		wait for 10 ns;
		t_blur_matrix_int <= (51,38,43,48,48,56,60,62,55,42,35,43,51,52,60,62,51,45,37,45,48,56,62,61,49,36,40,47,51,55,62,63,50,44,40,49,50,60,62,68,51,41,44,48,46,58,59,61,54,49,43,44,51,57,61,58,55,42,39,45,52,60,60,62);
		wait for 10 ns;
		t_blur_matrix_int <= (65,65,61,63,65,62,64,66,61,62,62,71,68,61,63,70,64,62,65,65,65,63,65,69,60,68,64,61,60,65,65,65,62,61,69,65,67,61,67,66,59,63,65,63,66,61,67,65,61,60,63,64,61,66,64,68,61,66,61,65,62,64,68,65);
		wait for 10 ns;
		t_blur_matrix_int <= (61,66,64,64,62,61,62,59,61,64,65,61,64,63,63,60,61,61,63,63,66,59,61,63,61,65,64,63,68,65,67,61,65,64,65,63,65,59,62,60,64,62,68,61,65,61,63,60,64,58,64,65,66,59,59,60,65,66,64,68,63,60,64,64);
		wait for 10 ns;
		t_blur_matrix_int <= (52,45,43,155,210,181,194,169,57,46,44,154,196,203,175,189,58,52,42,121,213,184,191,176,60,52,44,90,205,199,182,190,58,51,43,58,202,195,195,189,58,58,44,47,181,203,192,192,63,60,54,46,143,201,186,193,65,60,51,38,95,208,196,184);
		wait for 10 ns;
		t_blur_matrix_int <= (181,158,154,131,117,125,112,133,175,170,158,140,114,97,120,108,186,179,154,134,107,101,83,127,189,177,161,132,100,80,97,94,182,186,165,144,93,82,73,112,188,189,163,130,110,74,89,138,183,197,168,133,94,96,119,109,186,177,175,134,125,91,100,119);
		wait for 10 ns;
		t_blur_matrix_int <= (112,105,82,80,91,83,80,91,148,97,76,75,83,94,82,99,104,78,72,75,81,91,92,91,99,85,83,82,77,84,99,69,108,100,82,90,83,89,78,77,107,124,86,94,88,79,66,84,125,94,115,93,70,71,77,83,118,127,101,90,68,80,78,94);
		wait for 10 ns;
		t_blur_matrix_int <= (101,96,77,93,88,109,113,110,95,69,82,88,104,111,106,104,66,78,89,102,113,103,104,102,82,81,94,106,104,103,102,103,83,91,109,107,104,102,104,100,89,101,102,110,105,109,101,89,100,100,108,104,104,102,80,93,106,102,97,109,97,90,89,96);
		wait for 10 ns;
		t_blur_matrix_int <= (105,100,110,101,90,88,96,101,106,108,102,86,90,101,96,102,107,109,90,100,96,103,100,107,102,84,95,100,101,106,100,99,90,88,92,100,105,107,106,101,92,94,97,99,103,104,98,95,96,90,103,101,103,103,96,90,93,94,99,106,99,89,84,110);
		wait for 10 ns;
		t_blur_matrix_int <= (104,106,110,108,96,109,117,121,106,102,101,94,108,121,106,116,107,98,90,106,111,117,110,107,105,96,101,109,114,108,109,100,88,96,108,113,106,104,108,73,94,104,109,105,106,91,74,90,110,107,106,107,98,69,92,100,117,104,107,98,96,54,106,106);
		wait for 10 ns;
		t_blur_matrix_int <= (119,123,104,82,110,111,110,92,122,97,80,120,123,107,92,69,93,81,104,109,113,92,65,78,72,90,111,110,96,81,88,103,97,106,100,92,79,86,98,85,103,104,101,83,78,101,94,84,102,107,96,79,75,71,48,46,103,84,68,55,40,38,51,70);
		wait for 10 ns;
		t_blur_matrix_int <= (89,84,74,71,68,62,37,78,75,77,60,48,39,37,34,71,85,66,66,79,80,58,65,93,80,74,101,106,94,54,48,65,86,79,87,61,55,34,42,45,75,45,38,27,32,30,26,32,50,48,46,29,30,32,30,42,58,47,32,22,21,19,31,76);
		wait for 10 ns;
		t_blur_matrix_int <= (137,147,140,140,108,103,109,101,127,132,135,126,110,115,92,82,99,107,108,120,103,80,47,42,67,62,104,92,57,53,52,34,43,69,87,78,84,59,50,66,49,77,80,112,70,81,71,104,84,74,110,67,60,34,58,65,98,88,82,50,19,24,39,83);
		wait for 10 ns;
		t_blur_matrix_int <= (105,100,73,56,73,96,98,110,86,63,60,61,87,57,46,49,36,40,56,99,76,31,53,42,33,82,88,43,43,43,47,53,86,59,49,66,45,36,62,49,59,90,87,29,40,27,63,68,79,88,48,60,61,18,66,64,53,54,72,61,33,14,67,41);
		wait for 10 ns;
		t_blur_matrix_int <= (86,76,67,35,54,36,69,70,48,39,42,22,24,26,21,25,24,23,23,15,22,22,20,19,23,19,16,10,24,22,29,96,34,21,14,11,10,17,68,164,15,14,20,12,23,95,161,150,12,8,14,43,110,173,134,90,14,12,31,120,160,126,94,117);
		wait for 10 ns;
		t_blur_matrix_int <= (13,52,133,136,166,174,143,136,15,35,135,184,157,129,139,151,35,109,174,150,125,144,176,186,133,171,138,120,143,188,194,197,160,117,117,154,172,187,189,189,92,105,166,187,176,176,175,180,101,160,185,185,173,169,172,172,168,176,181,172,164,166,168,177);
		wait for 10 ns;
		t_blur_matrix_int <= (146,167,181,177,188,189,188,182,180,191,191,186,187,187,182,181,188,190,187,183,189,184,184,184,192,186,187,181,187,180,181,182,185,187,185,184,183,186,183,182,183,186,184,181,183,181,177,181,182,184,182,178,180,183,171,176,180,180,178,181,180,173,177,179);
		wait for 10 ns;
		t_blur_matrix_int <= (183,186,186,186,186,186,182,185,186,188,189,181,183,183,183,185,188,188,184,185,179,182,187,186,186,183,187,185,182,184,184,189,187,188,183,185,183,183,185,182,179,184,184,182,183,182,184,185,184,181,179,181,179,186,184,186,178,180,179,181,183,183,184,185);
		wait for 10 ns;
		t_blur_matrix_int <= (187,188,191,191,192,192,193,193,187,186,192,191,192,193,191,192,187,191,190,191,191,193,190,191,185,189,189,189,190,190,193,182,186,190,186,187,191,194,198,192,184,187,188,192,190,195,190,191,188,187,187,189,191,190,190,191,186,189,188,188,193,193,174,123);
		wait for 10 ns;
		t_blur_matrix_int <= (194,194,198,198,193,194,196,195,191,196,199,196,197,198,198,195,189,200,198,197,199,197,199,192,191,200,195,200,200,189,149,92,197,201,202,194,139,77,65,57,198,198,180,107,68,62,66,61,170,128,112,99,63,61,66,57,78,81,118,108,85,66,66,62);
		wait for 10 ns;
		t_blur_matrix_int <= (197,200,205,198,169,141,109,82,199,198,175,144,111,79,57,54,170,118,87,67,62,62,56,58,68,58,60,59,67,59,61,60,56,57,53,60,65,60,65,72,61,57,57,62,71,85,93,110,60,60,64,77,104,118,134,138,74,97,107,129,137,139,149,151);
		wait for 10 ns;
		t_blur_matrix_int <= (50,58,63,66,65,92,135,181,55,56,60,69,84,128,173,198,56,63,65,89,129,166,183,203,67,83,100,137,169,180,192,188,87,124,144,166,186,192,115,40,134,157,176,189,196,115,19,17,154,168,180,193,157,27,19,21,159,172,192,147,35,13,19,22);
		wait for 10 ns;
		t_blur_matrix_int <= (208,211,76,15,14,26,18,22,211,144,17,13,14,21,25,23,195,46,36,17,19,25,21,26,79,15,21,16,20,25,27,20,17,11,16,20,21,24,22,21,15,18,19,23,27,23,17,17,20,20,19,26,23,27,18,18,21,20,30,28,28,26,16,18);
		wait for 10 ns;
		t_blur_matrix_int <= (20,24,20,15,16,26,27,27,20,27,17,19,16,26,30,21,23,25,19,24,23,28,21,20,27,26,23,18,27,27,20,21,22,21,27,27,28,28,20,15,25,15,24,24,32,30,22,22,18,22,29,32,38,39,25,28,17,16,25,34,24,39,37,40);
		wait for 10 ns;
		t_blur_matrix_int <= (22,23,37,76,111,124,125,119,19,23,58,96,121,128,120,118,14,26,73,111,126,121,118,114,16,41,88,119,124,119,119,120,18,63,107,126,123,120,118,128,37,84,115,124,124,117,121,132,60,99,122,123,123,116,129,142,81,116,125,123,121,120,133,144);
		wait for 10 ns;
		t_blur_matrix_int <= (118,124,133,139,143,140,139,137,118,131,137,142,139,138,141,136,124,134,139,142,141,141,140,138,131,141,145,139,140,141,139,138,137,142,144,142,143,139,139,142,141,143,143,141,141,141,135,139,147,146,146,143,142,143,138,142,146,143,144,142,142,141,142,139);
		wait for 10 ns;
		t_blur_matrix_int <= (139,137,138,137,134,133,136,135,139,138,139,133,135,133,134,135,138,138,139,139,138,137,133,134,139,140,139,138,136,136,138,137,138,140,139,139,138,138,135,134,140,140,138,141,137,140,134,137,139,138,142,140,137,137,136,137,141,139,140,141,139,140,139,140);
		wait for 10 ns;
		t_blur_matrix_int <= (136,132,133,134,135,133,131,131,136,135,133,134,132,133,135,134,138,128,129,132,135,134,136,135,135,134,133,134,132,131,135,134,136,136,136,136,135,132,131,134,135,136,134,133,134,131,135,133,138,136,135,137,136,137,136,134,139,137,133,135,136,133,134,133);
		wait for 10 ns;
		t_blur_matrix_int <= (133,132,132,133,132,130,135,129,134,131,135,133,134,134,132,131,134,133,132,132,134,134,135,130,133,134,135,133,130,129,132,131,134,135,132,133,133,132,130,131,130,132,134,133,132,134,132,134,134,135,135,135,133,132,134,128,135,134,135,134,132,129,130,127);
		wait for 10 ns;
		t_blur_matrix_int <= (76,70,73,72,70,68,71,64,76,70,71,68,72,68,69,64,76,76,71,69,71,71,72,64,74,73,73,72,68,69,69,68,69,73,71,72,73,66,67,65,79,75,75,75,71,72,72,66,72,73,73,79,76,72,71,69,79,77,75,73,70,69,71,68);
		wait for 10 ns;
		t_blur_matrix_int <= (66,66,66,67,76,86,101,116,65,64,64,66,74,84,97,113,66,68,65,70,74,84,94,112,67,68,65,66,73,85,98,110,66,65,67,71,69,79,93,110,65,65,69,64,68,79,93,108,63,64,62,61,67,81,92,109,67,66,61,61,63,75,92,106);
		wait for 10 ns;
		t_blur_matrix_int <= (124,132,142,148,149,148,146,148,124,132,141,146,150,150,148,152,121,136,141,151,150,149,148,149,122,133,140,149,149,149,149,150,122,135,146,148,153,146,149,147,122,139,144,150,147,146,148,151,123,132,143,148,151,148,148,152,121,133,142,141,151,149,151,153);
		wait for 10 ns;
		t_blur_matrix_int <= (148,149,145,137,125,114,97,76,146,148,147,139,129,115,94,74,150,148,149,139,127,111,96,76,149,147,147,137,129,114,98,78,148,150,149,141,131,113,101,75,147,152,147,137,129,112,97,75,154,150,147,137,129,118,96,74,152,151,147,142,128,113,98,76);
		wait for 10 ns;
		t_blur_matrix_int <= (55,43,43,48,50,53,57,59,56,42,41,45,49,53,58,61,56,41,40,46,55,53,59,63,55,41,42,46,54,59,60,62,54,36,36,43,47,57,55,60,51,40,38,46,52,54,58,62,51,43,40,47,53,47,56,60,50,41,40,45,46,53,58,60);
		wait for 10 ns;
		t_blur_matrix_int <= (61,61,63,63,64,60,64,63,64,63,59,65,67,65,64,65,61,62,61,64,66,65,68,65,61,61,62,64,62,64,65,64,63,62,58,60,62,60,68,67,62,59,63,60,62,60,59,59,59,61,63,66,64,65,60,61,55,66,62,65,63,62,61,65);
		wait for 10 ns;
		t_blur_matrix_int <= (67,62,67,65,69,62,66,65,65,64,66,61,60,60,64,66,67,66,63,66,64,61,65,66,61,61,62,65,65,63,68,68,61,62,62,62,63,62,69,67,63,65,59,64,64,63,70,67,62,62,60,62,64,66,68,70,65,63,62,62,67,68,67,70);
		wait for 10 ns;
		t_blur_matrix_int <= (65,61,58,45,55,193,197,189,65,67,59,47,43,142,204,187,66,65,59,52,45,111,210,191,68,69,64,57,47,70,192,198,70,67,67,62,57,52,118,216,69,72,69,67,60,52,65,182,71,71,73,67,67,57,51,97,73,71,70,71,67,64,55,53);
		wait for 10 ns;
		t_blur_matrix_int <= (175,189,172,164,125,108,92,127,186,173,189,159,156,132,113,104,179,193,175,187,152,135,153,114,199,177,195,162,136,161,144,139,193,205,180,160,135,157,160,142,211,194,199,166,132,153,159,156,197,208,197,174,167,152,167,165,149,208,195,177,183,170,173,125);
		wait for 10 ns;
		t_blur_matrix_int <= (103,121,104,71,69,85,94,110,127,91,91,76,80,83,104,104,141,94,64,80,96,100,106,103,108,92,65,91,90,95,104,106,95,55,80,98,100,90,96,101,101,66,93,104,100,98,93,90,103,99,95,98,100,100,90,82,61,121,93,85,97,98,90,85);
		wait for 10 ns;
		t_blur_matrix_int <= (101,104,105,101,79,87,92,97,106,99,96,75,75,92,93,98,107,100,73,70,85,91,95,94,99,88,80,95,91,94,96,90,81,67,99,96,92,98,86,89,79,83,91,93,97,91,89,88,83,92,98,101,96,96,89,92,88,95,100,94,110,102,96,96);
		wait for 10 ns;
		t_blur_matrix_int <= (94,93,95,101,95,89,95,106,99,101,90,93,87,85,109,105,91,95,93,85,88,107,99,76,88,99,91,84,103,108,106,104,85,90,86,100,102,110,107,106,91,90,92,108,99,93,85,77,85,92,106,97,82,82,83,87,86,91,94,98,96,94,85,66);
		wait for 10 ns;
		t_blur_matrix_int <= (102,107,106,106,104,63,104,101,101,99,104,114,110,69,97,83,65,70,96,111,106,69,65,42,91,74,58,69,86,70,38,37,71,45,70,54,42,58,57,43,64,37,33,33,52,54,38,62,74,72,60,58,37,35,53,65,61,58,52,45,45,58,73,63);
		wait for 10 ns;
		t_blur_matrix_int <= (77,62,43,27,33,74,76,39,47,36,27,50,76,55,25,23,48,36,56,65,35,36,19,18,45,59,47,42,34,31,24,36,51,63,50,41,31,22,38,79,59,46,37,31,16,22,82,60,36,26,20,13,23,50,103,49,32,22,15,12,22,60,102,31);
		wait for 10 ns;
		t_blur_matrix_int <= (31,28,29,18,30,17,59,105,19,30,24,18,23,22,87,86,34,34,12,18,21,60,106,46,46,16,11,16,41,73,72,25,25,11,11,25,62,58,50,19,14,13,15,40,71,49,25,16,11,13,17,42,73,47,16,26,14,18,25,41,45,46,22,23);
		wait for 10 ns;
		t_blur_matrix_int <= (93,89,50,20,13,24,91,69,79,49,22,25,24,86,92,41,51,26,17,33,86,101,68,64,29,27,25,70,80,51,93,93,22,23,35,78,42,67,79,49,23,38,40,44,26,45,80,19,30,23,29,22,20,63,71,11,35,23,26,21,17,70,60,15);
		wait for 10 ns;
		t_blur_matrix_int <= (44,73,76,21,14,14,86,64,59,64,28,11,23,17,91,50,81,19,15,52,8,29,87,75,37,14,70,67,4,54,124,153,13,61,120,22,14,105,147,123,18,127,97,9,47,135,93,92,31,125,54,75,105,81,79,104,72,107,95,127,108,54,97,145);
		wait for 10 ns;
		t_blur_matrix_int <= (16,47,126,158,113,102,133,179,60,141,151,107,96,137,177,188,138,144,99,104,147,172,186,188,121,95,99,148,183,179,185,184,89,102,152,183,189,184,179,179,108,164,180,186,186,182,180,179,170,183,187,182,182,183,175,174,177,180,182,181,183,180,171,173);
		wait for 10 ns;
		t_blur_matrix_int <= (183,181,175,169,166,168,176,175,182,174,175,167,165,170,174,171,173,170,166,164,168,175,171,172,173,166,165,167,169,170,173,167,175,170,166,169,170,163,170,170,178,170,172,169,167,172,173,161,171,170,167,164,171,169,172,163,170,164,168,167,168,171,165,158);
		wait for 10 ns;
		t_blur_matrix_int <= (176,174,178,177,177,174,174,174,171,172,169,177,172,170,175,176,167,166,170,166,168,172,172,174,171,166,166,169,158,167,178,180,164,160,163,165,164,165,174,180,163,157,162,168,169,167,175,182,151,154,167,170,167,169,176,178,159,161,171,174,171,171,177,174);
		wait for 10 ns;
		t_blur_matrix_int <= (179,181,182,178,180,182,185,186,176,178,180,181,182,184,183,188,177,182,184,180,181,185,187,186,179,179,176,180,184,185,184,183,180,186,182,178,182,182,168,102,183,180,180,178,173,166,146,89,176,179,170,165,175,177,162,129,170,166,164,175,176,179,171,144);
		wait for 10 ns;
		t_blur_matrix_int <= (185,190,193,189,185,139,70,65,190,193,189,142,61,60,71,61,187,163,73,60,24,59,108,83,130,30,30,75,64,43,119,107,45,25,25,70,86,56,75,124,49,56,60,45,75,82,68,96,65,45,56,80,60,67,70,67,93,61,50,51,98,82,77,83);
		wait for 10 ns;
		t_blur_matrix_int <= (87,86,116,120,108,96,103,109,85,78,105,120,127,138,136,137,84,82,96,124,134,143,138,142,84,100,81,115,134,137,136,146,92,108,93,103,129,123,135,147,117,93,104,82,123,129,130,142,115,102,97,76,107,127,128,148,95,123,101,100,106,128,137,164);
		wait for 10 ns;
		t_blur_matrix_int <= (127,139,143,146,147,143,141,154,143,141,144,140,150,146,154,168,143,145,142,144,152,159,177,197,148,146,151,155,165,178,191,169,147,151,157,161,178,188,113,38,146,149,162,186,180,83,15,16,159,173,186,163,55,19,17,19,180,182,117,42,20,19,14,19);
		wait for 10 ns;
		t_blur_matrix_int <= (166,191,145,27,16,18,18,20,195,162,32,14,13,16,20,26,163,40,16,14,11,21,24,23,41,16,18,16,21,20,23,25,21,11,14,16,18,23,26,24,19,9,19,19,21,20,20,31,16,14,20,22,27,25,22,29,16,18,22,29,28,25,22,28);
		wait for 10 ns;
		t_blur_matrix_int <= (22,31,29,23,30,23,26,20,32,32,26,24,24,17,25,21,25,31,29,30,31,21,18,19,29,27,25,26,26,22,18,24,26,31,31,32,21,23,20,18,32,33,37,27,24,24,18,18,28,32,26,21,18,23,18,17,28,26,29,21,21,23,17,22);
		wait for 10 ns;
		t_blur_matrix_int <= (14,16,29,32,34,27,25,50,24,23,29,23,14,23,28,79,21,26,28,30,20,29,42,93,22,25,25,25,26,27,65,106,22,24,23,25,26,40,80,111,23,28,26,22,34,52,93,114,29,29,24,37,40,71,104,110,29,25,27,35,52,87,112,110);
		wait for 10 ns;
		t_blur_matrix_int <= (99,120,123,124,113,121,140,146,110,124,121,121,116,127,146,147,123,122,119,120,122,137,147,144,121,120,116,118,130,143,144,147,118,120,110,121,137,146,148,148,110,112,107,126,143,147,149,148,107,106,111,134,150,151,146,148,102,99,118,141,148,150,150,149);
		wait for 10 ns;
		t_blur_matrix_int <= (144,147,143,147,147,145,144,142,143,146,147,148,147,145,142,140,149,144,145,147,147,145,143,141,149,146,145,149,148,145,146,142,144,151,144,143,146,147,146,144,149,147,147,150,145,141,144,145,146,145,144,144,143,142,142,143,147,142,142,145,145,141,143,144);
		wait for 10 ns;
		t_blur_matrix_int <= (143,143,141,140,140,138,135,137,142,140,140,140,138,142,136,139,143,142,141,138,137,138,137,138,142,146,144,141,142,140,140,138,144,143,144,142,138,139,136,139,146,142,143,143,140,141,139,139,144,144,144,142,140,140,143,140,146,145,142,144,141,139,140,141);
		wait for 10 ns;
		t_blur_matrix_int <= (138,134,134,134,136,135,135,134,137,136,135,133,137,135,133,135,138,139,135,137,135,135,135,137,137,133,136,136,138,137,136,136,138,139,136,138,138,135,135,137,137,137,139,134,138,138,135,136,140,141,141,139,138,140,137,137,137,135,139,143,141,140,135,137);
		wait for 10 ns;
		t_blur_matrix_int <= (135,136,136,135,134,131,130,130,134,139,135,133,135,131,130,129,133,133,133,132,133,131,131,129,136,133,133,132,136,133,133,130,135,136,135,132,136,130,132,129,137,134,133,130,133,130,131,131,137,136,135,134,135,131,126,129,136,138,133,138,134,133,135,132);
		wait for 10 ns;
		t_blur_matrix_int <= (75,74,76,75,70,72,69,67,75,76,78,75,71,65,70,71,72,77,75,70,70,72,68,65,72,75,72,70,72,70,69,66,75,71,72,73,70,74,72,62,74,76,68,75,74,74,71,69,72,73,74,74,74,69,70,67,67,71,73,70,72,67,68,66);
		wait for 10 ns;
		t_blur_matrix_int <= (63,68,62,59,63,72,92,107,68,63,61,58,57,74,93,107,66,63,61,59,59,74,91,105,65,65,62,54,58,73,88,106,64,63,58,55,60,76,90,104,65,66,58,58,55,70,91,104,64,65,63,59,59,73,90,105,69,69,63,55,62,73,90,105);
		wait for 10 ns;
		t_blur_matrix_int <= (117,135,146,149,150,150,150,148,122,135,140,151,153,148,151,153,122,130,141,146,151,153,151,150,118,128,143,145,149,146,148,151,116,129,140,148,153,149,152,155,117,130,140,145,147,152,152,152,119,129,139,146,148,150,150,152,120,130,141,146,152,149,148,154);
		wait for 10 ns;
		t_blur_matrix_int <= (154,154,148,141,128,116,96,75,151,151,149,141,128,118,101,75,152,153,148,143,129,114,99,79,154,150,152,142,130,115,98,76,152,153,151,141,128,117,102,79,152,152,148,139,128,116,95,77,150,148,148,139,131,115,101,79,151,151,148,140,131,123,99,79);
		wait for 10 ns;
		t_blur_matrix_int <= (55,42,39,44,48,52,55,61,53,38,35,43,50,51,57,56,55,37,38,41,49,50,57,53,51,38,38,48,44,48,60,58,51,40,37,45,51,56,61,56,50,41,41,37,53,54,61,59,59,44,37,43,49,51,63,59,60,42,34,45,48,52,60,58);
		wait for 10 ns;
		t_blur_matrix_int <= (58,67,64,62,62,61,63,64,58,63,60,62,64,60,62,63,62,61,63,61,62,63,62,58,59,65,65,64,66,65,65,64,64,63,63,63,67,70,66,65,64,65,62,65,67,64,62,67,62,64,67,65,65,68,67,64,62,63,65,65,64,64,68,66);
		wait for 10 ns;
		t_blur_matrix_int <= (59,65,66,67,65,69,68,70,65,64,62,63,64,68,68,72,61,63,63,64,64,65,68,71,63,65,62,64,67,67,70,68,62,62,60,61,64,65,70,71,64,63,65,63,65,68,69,73,64,63,66,65,69,72,69,73,63,65,64,66,69,68,68,74);
		wait for 10 ns;
		t_blur_matrix_int <= (73,72,76,74,74,69,55,52,74,75,79,75,75,69,66,55,69,75,81,77,74,71,66,58,77,79,76,74,77,73,69,58,74,78,76,80,76,71,67,61,77,80,84,79,78,74,74,61,74,76,76,79,78,74,74,64,73,76,83,84,77,76,74,67);
		wait for 10 ns;
		t_blur_matrix_int <= (77,199,189,183,179,176,182,102,55,167,217,192,180,180,186,119,54,151,209,210,192,186,180,155,50,149,211,205,200,188,181,134,51,145,212,204,208,200,168,82,52,139,210,208,202,202,125,69,56,113,214,208,205,185,87,68,62,80,200,209,211,155,70,74);
		wait for 10 ns;
		t_blur_matrix_int <= (103,111,84,80,92,87,78,96,116,93,89,83,86,71,76,89,104,87,93,93,74,68,82,96,87,89,90,92,84,82,92,92,70,89,94,86,85,92,91,88,66,84,86,84,89,91,93,73,69,74,82,80,83,83,74,81,75,76,75,85,82,85,88,96);
		wait for 10 ns;
		t_blur_matrix_int <= (95,96,101,93,93,89,82,93,97,99,94,77,82,73,93,97,94,93,87,84,81,103,102,98,84,84,82,96,108,103,96,92,70,78,96,106,100,98,99,96,77,93,103,99,101,99,85,87,92,91,90,78,101,85,81,92,91,97,97,65,81,78,81,70);
		wait for 10 ns;
		t_blur_matrix_int <= (100,93,86,81,95,81,65,49,95,93,98,105,88,69,37,36,91,69,73,103,91,68,41,44,91,72,78,83,63,53,45,44,80,59,50,54,29,35,65,45,94,42,17,27,20,45,52,26,92,59,18,15,28,61,32,21,67,55,16,18,54,64,18,16);
		wait for 10 ns;
		t_blur_matrix_int <= (37,54,44,58,58,68,73,44,46,38,48,47,58,69,59,47,42,29,33,32,49,65,55,42,35,28,21,21,43,52,46,39,24,22,21,19,27,55,42,48,17,22,23,22,23,55,62,36,21,17,19,23,20,34,56,46,13,25,22,24,21,25,33,56);
		wait for 10 ns;
		t_blur_matrix_int <= (27,28,21,14,26,77,85,21,34,30,25,18,35,54,65,33,32,22,25,28,45,35,53,62,51,40,33,23,51,19,56,84,58,62,30,24,51,20,34,81,50,65,32,20,53,29,15,61,37,56,45,21,57,31,12,24,41,42,44,33,61,39,26,30);
		wait for 10 ns;
		t_blur_matrix_int <= (15,25,69,21,26,25,28,33,32,39,51,17,22,22,24,31,62,34,20,22,19,18,20,22,76,36,14,20,26,20,22,22,104,58,17,21,20,24,21,15,97,105,38,24,19,21,18,17,66,119,72,66,68,30,11,14,45,127,40,25,32,21,15,10);
		wait for 10 ns;
		t_blur_matrix_int <= (57,61,61,61,36,88,55,41,25,34,36,26,24,63,40,43,27,22,20,16,13,43,43,69,31,19,21,16,18,53,81,76,22,19,9,13,38,78,94,48,11,8,14,33,100,88,75,63,10,12,28,107,125,69,73,129,6,21,108,127,83,84,136,165);
		wait for 10 ns;
		t_blur_matrix_int <= (82,80,95,109,93,96,156,158,64,65,76,122,94,154,143,162,59,46,75,93,109,125,137,160,59,55,111,126,146,152,155,163,66,97,134,122,165,168,163,168,128,135,130,137,171,166,167,172,157,132,107,141,177,163,169,179,141,140,108,130,171,163,156,181);
		wait for 10 ns;
		t_blur_matrix_int <= (176,175,174,175,180,176,172,169,169,164,164,172,177,170,164,157,165,157,165,168,170,162,158,154,162,166,175,174,166,156,152,151,170,176,177,169,162,151,145,151,178,178,175,167,151,146,140,148,182,183,168,155,148,144,141,147,175,172,161,152,146,145,143,151);
		wait for 10 ns;
		t_blur_matrix_int <= (167,166,167,164,167,161,160,162,158,159,165,157,158,161,164,163,150,167,158,159,162,162,161,160,159,161,163,166,166,156,154,163,154,155,166,167,159,144,146,155,152,159,171,163,153,136,146,154,156,169,170,157,142,141,150,151,166,173,153,130,136,145,150,159);
		wait for 10 ns;
		t_blur_matrix_int <= (161,160,171,172,172,170,173,169,162,159,165,164,167,170,177,178,161,164,154,163,175,181,183,175,161,151,160,174,176,180,186,179,151,163,173,182,179,186,190,182,163,169,174,179,182,183,188,184,166,168,175,183,177,183,189,186,168,173,177,182,180,185,189,189);
		wait for 10 ns;
		t_blur_matrix_int <= (173,169,175,180,185,185,174,159,177,176,180,180,182,188,182,175,178,176,181,181,179,181,181,179,182,180,184,181,183,183,186,178,181,179,182,182,186,182,182,177,184,181,183,184,188,188,186,184,186,186,188,190,192,192,190,190,186,188,189,192,199,197,197,196);
		wait for 10 ns;
		t_blur_matrix_int <= (113,72,58,54,60,108,75,63,139,93,59,55,46,43,97,58,155,110,69,54,45,31,48,78,157,119,76,60,45,34,14,52,157,134,88,57,44,33,19,21,167,139,89,59,49,27,19,17,176,147,109,65,56,30,13,19,182,160,123,73,55,38,13,17);
		wait for 10 ns;
		t_blur_matrix_int <= (57,111,113,112,106,123,148,168,56,66,118,113,112,125,138,114,64,38,102,110,119,124,128,103,70,46,65,111,112,129,132,111,72,52,53,107,110,117,127,116,33,56,44,93,120,129,130,121,20,57,41,70,131,129,143,117,20,37,46,50,125,134,149,113);
		wait for 10 ns;
		t_blur_matrix_int <= (144,72,26,16,18,20,20,19,88,41,13,12,14,23,18,21,80,40,13,13,19,15,17,18,77,26,20,15,11,14,19,17,71,24,19,15,17,21,21,20,46,23,27,25,19,22,20,18,37,19,18,21,17,21,21,23,31,18,22,15,23,20,19,25);
		wait for 10 ns;
		t_blur_matrix_int <= (13,20,28,29,33,27,27,30,22,21,24,29,29,30,31,32,26,26,26,30,30,31,29,28,29,32,29,26,30,31,37,36,22,31,27,32,28,30,35,30,26,24,33,31,31,44,33,37,22,27,30,28,36,34,36,30,27,30,29,31,31,40,38,26);
		wait for 10 ns;
		t_blur_matrix_int <= (27,29,27,17,14,20,18,24,29,32,23,15,20,22,24,24,29,23,21,15,14,23,28,26,28,21,21,16,17,19,24,22,28,22,26,18,15,20,27,23,26,21,17,19,20,22,20,17,21,19,21,15,20,25,21,26,19,16,18,20,22,25,16,23);
		wait for 10 ns;
		t_blur_matrix_int <= (30,23,34,41,63,100,112,104,24,21,32,47,78,106,112,102,22,27,39,60,101,112,107,97,23,29,43,78,102,112,105,97,20,24,60,97,114,112,106,101,24,31,73,106,119,112,101,106,26,48,92,117,117,110,106,121,33,65,105,119,113,106,111,130);
		wait for 10 ns;
		t_blur_matrix_int <= (99,106,127,147,149,151,151,147,105,109,135,148,154,148,151,149,101,115,136,149,148,148,151,147,105,127,137,146,149,150,149,146,115,134,140,145,143,149,146,147,125,134,133,133,144,148,148,147,130,133,128,131,134,137,144,146,135,133,131,128,132,131,134,137);
		wait for 10 ns;
		t_blur_matrix_int <= (143,143,145,147,145,144,146,146,147,144,147,145,141,148,144,144,147,146,151,144,145,144,146,147,148,149,146,143,146,143,145,144,145,146,145,147,140,143,144,143,146,150,147,145,144,140,139,142,149,149,147,148,145,143,145,142,138,142,146,142,143,143,144,141);
		wait for 10 ns;
		t_blur_matrix_int <= (140,142,142,144,140,141,140,139,144,142,141,145,143,144,142,140,146,143,142,144,143,142,141,145,145,146,143,141,143,143,138,140,144,141,145,147,143,143,143,142,143,143,143,144,143,145,142,141,142,141,140,144,145,146,142,141,139,141,141,144,143,146,143,140);
		wait for 10 ns;
		t_blur_matrix_int <= (141,139,140,138,139,136,138,136,143,143,142,139,138,139,138,137,143,144,142,139,137,137,137,138,140,142,142,138,143,135,138,139,144,139,138,142,138,139,142,139,140,139,142,138,137,136,139,137,141,138,140,138,136,139,140,138,141,140,139,140,134,137,136,137);
		wait for 10 ns;
		t_blur_matrix_int <= (138,136,136,133,135,131,132,128,136,136,138,131,134,131,128,132,136,137,135,133,137,131,131,130,138,138,138,135,133,132,135,128,135,138,136,134,135,130,126,128,136,140,136,134,134,133,133,126,136,139,135,135,134,133,131,126,139,140,136,136,134,132,130,127);
		wait for 10 ns;
		t_blur_matrix_int <= (69,72,70,72,71,71,69,69,65,73,72,67,72,70,68,67,73,76,73,75,70,68,68,69,68,72,73,70,69,62,67,66,72,75,71,72,69,62,63,69,69,72,71,70,68,66,65,65,67,72,68,67,68,67,65,62,67,71,66,72,69,68,68,60);
		wait for 10 ns;
		t_blur_matrix_int <= (64,67,63,57,59,73,91,106,68,65,62,59,61,71,88,106,66,70,62,57,59,74,89,106,66,64,58,57,66,71,87,105,63,62,60,57,60,71,88,100,61,61,59,54,51,70,89,102,66,64,60,54,57,70,89,104,64,68,61,55,58,68,89,103);
		wait for 10 ns;
		t_blur_matrix_int <= (119,131,138,144,148,151,149,151,118,133,139,149,149,150,152,152,115,131,141,148,151,150,152,152,116,129,140,148,148,153,155,153,115,129,140,145,151,151,155,156,118,130,141,149,152,153,152,157,118,122,139,147,151,154,155,153,117,127,143,151,152,153,155,154);
		wait for 10 ns;
		t_blur_matrix_int <= (155,150,152,144,131,117,102,81,155,152,150,146,130,117,100,79,151,153,150,145,132,116,100,80,151,154,154,143,130,117,102,84,153,153,151,145,130,116,103,80,154,153,149,143,131,115,103,78,154,151,150,139,134,122,103,78,157,158,151,144,132,116,101,78);
		wait for 10 ns;
		t_blur_matrix_int <= (56,43,41,45,46,52,62,60,60,44,41,42,48,48,57,59,63,45,40,46,49,54,60,66,62,49,45,51,52,55,64,64,60,46,47,52,59,61,63,59,58,43,45,45,60,57,62,62,56,47,42,47,56,57,64,61,58,43,43,48,51,54,61,64);
		wait for 10 ns;
		t_blur_matrix_int <= (62,67,67,67,66,68,68,64,64,66,71,68,68,73,68,71,67,67,65,71,73,73,67,69,68,66,67,67,70,65,68,66,64,65,70,68,68,68,67,67,64,66,69,66,68,67,71,70,68,70,66,65,69,70,73,68,69,64,70,66,72,70,71,71);
		wait for 10 ns;
		t_blur_matrix_int <= (68,67,66,66,68,67,63,70,64,63,66,64,64,62,71,118,68,63,64,64,67,63,88,111,65,63,65,68,68,72,80,80,68,69,68,67,71,68,77,92,69,69,70,66,69,70,74,94,66,67,67,66,70,74,73,80,70,65,66,69,72,71,74,78);
		wait for 10 ns;
		t_blur_matrix_int <= (109,81,79,81,78,79,75,73,131,73,77,83,79,79,76,74,80,79,82,79,81,78,82,81,78,81,80,84,80,86,80,81,77,77,80,87,83,82,85,82,77,85,79,84,85,84,86,88,82,80,78,80,81,80,81,82,82,82,82,79,79,78,76,75);
		wait for 10 ns;
		t_blur_matrix_int <= (62,62,171,213,212,129,80,76,70,67,116,221,210,110,79,78,76,72,84,185,215,126,76,81,81,76,70,123,221,155,84,83,82,78,76,86,188,172,88,87,84,81,79,82,125,161,89,83,79,81,91,98,89,113,75,83,75,80,108,86,56,78,84,70);
		wait for 10 ns;
		t_blur_matrix_int <= (82,83,78,80,70,75,103,97,88,87,82,64,75,102,95,94,80,81,84,77,92,87,96,94,77,71,86,92,92,94,84,104,79,71,101,90,92,98,100,90,70,94,98,102,95,97,104,99,84,98,106,102,104,99,95,82,99,89,100,101,94,102,93,72);
		wait for 10 ns;
		t_blur_matrix_int <= (87,84,83,54,47,57,49,36,103,84,70,65,50,53,48,22,101,99,81,75,70,56,29,23,93,85,68,66,32,24,25,36,92,59,62,40,26,26,47,60,77,53,23,24,23,32,74,52,57,26,29,45,14,12,70,33,45,16,49,41,12,11,81,39);
		wait for 10 ns;
		t_blur_matrix_int <= (46,51,28,20,68,47,18,17,33,33,17,23,82,37,19,18,26,16,15,28,79,25,14,19,27,13,17,14,74,30,23,27,17,16,15,15,54,55,41,33,11,19,18,13,29,72,31,18,13,45,22,19,11,29,50,24,26,44,16,27,16,18,31,74);
		wait for 10 ns;
		t_blur_matrix_int <= (15,33,21,33,21,24,21,40,28,40,30,30,20,22,31,21,47,32,27,27,19,26,30,18,29,24,38,19,24,30,29,26,26,35,33,19,26,28,21,29,27,59,32,20,24,22,18,41,58,50,21,14,24,23,14,55,70,31,15,14,29,14,19,69);
		wait for 10 ns;
		t_blur_matrix_int <= (46,34,34,39,60,35,44,27,31,37,28,29,65,67,74,27,24,37,26,22,52,81,98,49,34,28,14,36,62,64,50,70,48,30,13,23,75,45,45,41,38,36,17,21,46,22,54,24,23,51,22,18,21,31,72,28,14,30,46,26,25,22,100,37);
		wait for 10 ns;
		t_blur_matrix_int <= (36,117,45,16,12,12,9,7,20,85,75,15,13,10,11,13,24,53,103,16,8,9,13,68,58,67,141,50,7,11,53,128,18,29,124,42,7,38,118,113,9,9,81,82,26,110,118,84,8,4,28,84,99,130,89,90,7,6,15,69,111,84,83,140);
		wait for 10 ns;
		t_blur_matrix_int <= (15,91,142,84,83,136,171,148,78,136,98,79,131,161,154,147,137,104,88,125,168,153,166,155,104,87,114,171,150,162,169,165,84,101,160,150,151,163,175,173,100,151,139,143,157,161,178,173,141,144,139,138,145,164,177,172,158,134,137,138,142,155,176,177);
		wait for 10 ns;
		t_blur_matrix_int <= (143,141,118,131,155,149,155,180,145,148,121,140,166,150,168,182,147,152,127,139,155,161,171,182,161,164,134,135,148,153,175,190,165,166,130,124,147,158,180,188,175,168,134,109,158,174,184,170,177,172,148,108,159,178,171,153,172,174,163,134,167,168,148,148);
		wait for 10 ns;
		t_blur_matrix_int <= (164,168,155,154,155,149,148,155,180,166,150,153,155,157,155,156,182,162,151,155,155,151,146,125,184,153,153,152,144,141,122,124,166,149,143,147,145,122,128,129,153,140,138,141,124,128,134,133,141,133,127,127,126,132,135,138,135,127,134,139,135,133,139,139);
		wait for 10 ns;
		t_blur_matrix_int <= (165,137,122,136,142,150,157,166,133,121,137,141,145,151,160,170,122,126,139,145,146,155,164,175,130,133,143,146,145,155,165,171,137,143,147,150,148,155,166,170,143,147,150,150,153,154,160,166,145,149,145,153,152,156,160,166,146,150,149,151,154,159,156,163);
		wait for 10 ns;
		t_blur_matrix_int <= (168,177,178,187,182,188,188,188,166,176,179,183,183,187,185,188,174,175,180,187,184,183,189,189,177,176,178,181,186,186,191,192,177,180,180,181,186,186,190,189,177,177,176,182,184,184,192,189,175,178,180,182,186,184,184,187,173,175,180,182,181,180,182,181);
		wait for 10 ns;
		t_blur_matrix_int <= (187,186,189,194,195,199,199,199,186,191,195,197,195,197,197,200,187,190,197,195,198,198,201,199,190,188,194,196,198,197,199,200,191,192,194,195,197,199,201,199,190,190,194,197,199,196,201,202,189,189,192,196,196,198,200,200,187,187,191,189,194,196,198,199);
		wait for 10 ns;
		t_blur_matrix_int <= (191,171,134,84,61,41,17,11,191,176,147,97,64,43,23,21,190,181,155,110,68,45,25,16,197,185,163,122,72,51,32,16,200,193,173,127,84,59,36,20,203,195,178,138,97,60,45,26,201,199,186,150,106,66,58,38,200,193,189,165,116,72,56,38);
		wait for 10 ns;
		t_blur_matrix_int <= (15,25,45,38,102,138,155,122,13,12,30,43,68,133,150,129,7,11,21,52,44,139,147,130,13,11,18,47,37,138,147,128,15,17,18,30,44,106,150,132,20,16,14,23,52,78,151,149,22,16,14,16,59,61,149,152,20,12,16,18,45,50,138,155);
		wait for 10 ns;
		t_blur_matrix_int <= (33,26,26,23,24,27,34,28,55,29,31,19,24,22,23,31,64,29,27,37,24,27,25,29,65,31,26,26,27,31,26,26,75,35,22,22,24,31,30,29,76,25,22,20,27,30,29,38,70,32,36,17,28,33,32,34,89,37,28,21,25,30,28,29);
		wait for 10 ns;
		t_blur_matrix_int <= (28,27,30,32,41,36,32,23,33,28,35,33,39,39,29,25,30,34,33,35,42,34,26,22,36,32,33,37,40,37,29,18,32,35,30,34,40,33,31,21,36,29,33,35,31,27,28,23,33,37,37,40,34,22,24,25,33,40,40,36,32,25,18,23);
		wait for 10 ns;
		t_blur_matrix_int <= (20,22,21,25,29,28,17,20,20,17,22,26,27,25,16,19,17,20,23,27,29,23,18,26,21,22,23,26,25,19,19,42,22,25,26,32,28,19,24,66,20,22,29,24,19,18,28,77,28,26,30,21,16,28,62,99,24,26,28,20,18,29,77,107);
		wait for 10 ns;
		t_blur_matrix_int <= (39,85,117,122,109,100,123,136,50,98,120,114,108,112,130,142,67,108,120,115,103,121,137,149,91,118,120,112,107,124,142,148,108,121,117,110,113,132,148,147,115,122,115,109,123,141,149,149,118,117,110,112,124,146,147,145,119,113,110,114,131,144,146,146);
		wait for 10 ns;
		t_blur_matrix_int <= (142,133,134,130,131,130,129,130,140,137,132,132,132,128,129,128,144,139,138,136,133,133,134,131,146,144,139,137,137,132,131,130,146,147,146,145,144,138,137,136,145,146,145,142,144,143,143,142,143,143,144,146,143,142,150,148,142,141,142,141,141,143,145,148);
		wait for 10 ns;
		t_blur_matrix_int <= (132,132,135,139,142,139,140,144,128,130,127,128,133,132,139,139,133,128,129,129,134,130,132,130,130,128,125,128,127,130,130,129,133,135,134,131,133,132,130,128,141,136,135,134,133,134,134,129,141,144,144,141,140,134,136,137,148,144,147,148,141,138,135,136);
		wait for 10 ns;
		t_blur_matrix_int <= (143,140,142,144,145,144,145,140,138,140,140,140,140,140,143,144,132,131,136,140,139,143,142,141,126,125,129,130,131,137,139,141,125,127,127,127,124,126,133,131,127,128,126,127,130,129,127,126,132,128,124,125,129,130,125,126,133,132,126,128,130,131,125,125);
		wait for 10 ns;
		t_blur_matrix_int <= (141,141,140,143,135,139,137,136,143,139,140,137,141,136,136,136,142,142,140,139,136,138,135,137,139,141,138,135,136,137,135,134,134,134,138,137,131,133,131,133,129,127,125,130,131,131,133,130,122,124,125,122,124,126,126,132,125,125,121,119,120,122,126,124);
		wait for 10 ns;
		t_blur_matrix_int <= (137,136,135,133,134,129,130,127,135,135,134,133,134,133,129,128,135,135,131,133,132,129,128,123,134,131,134,132,130,126,128,124,132,134,134,136,131,130,129,124,134,128,133,131,131,130,127,125,129,132,133,137,130,131,127,127,124,132,134,129,130,129,129,128);
		wait for 10 ns;
		t_blur_matrix_int <= (67,72,69,69,67,62,67,60,63,72,65,65,67,64,67,63,71,68,69,68,64,66,64,64,63,67,65,66,68,67,64,66,64,71,68,66,68,67,68,63,71,70,68,68,72,66,67,68,66,66,72,66,73,74,69,70,65,69,69,70,75,70,71,65);
		wait for 10 ns;
		t_blur_matrix_int <= (63,66,62,53,57,68,88,105,60,63,59,56,57,70,86,108,62,65,61,59,56,68,85,105,68,63,59,59,60,67,88,102,66,64,60,61,54,65,87,105,68,64,60,60,56,66,83,102,65,63,65,53,55,64,84,97,67,62,57,54,51,67,86,103);
		wait for 10 ns;
		t_blur_matrix_int <= (123,134,142,147,148,152,156,154,118,130,140,147,149,151,152,155,113,131,139,148,151,152,154,155,119,130,140,144,153,153,156,156,120,129,140,146,151,152,156,156,117,128,140,150,152,149,155,154,117,122,137,147,155,148,153,154,118,129,137,150,154,151,153,154);
		wait for 10 ns;
		t_blur_matrix_int <= (155,154,151,146,131,115,98,75,156,155,155,145,131,119,102,78,154,155,151,144,133,117,100,77,154,156,150,146,132,121,99,80,157,155,154,144,135,122,104,77,156,157,153,145,130,119,104,81,155,155,156,147,133,120,102,82,154,157,158,147,136,124,109,83);
		wait for 10 ns;
		t_blur_matrix_int <= (59,46,39,46,53,53,61,62,57,47,41,45,51,58,59,63,58,47,40,49,53,55,61,63,57,48,43,50,54,49,57,62,53,44,43,48,54,52,65,59,57,44,47,50,55,57,56,62,58,44,50,48,56,58,65,62,57,44,41,51,50,55,62,65);
		wait for 10 ns;
		t_blur_matrix_int <= (66,68,70,64,70,67,69,69,69,66,66,69,72,69,68,66,65,71,69,69,69,62,69,66,64,64,70,70,71,71,67,67,64,68,71,69,66,67,74,70,63,67,75,68,70,65,64,64,64,74,70,66,68,65,66,64,68,68,68,65,68,65,68,66);
		wait for 10 ns;
		t_blur_matrix_int <= (68,70,68,67,72,74,75,75,67,69,66,64,71,71,76,79,67,66,66,71,71,73,76,80,67,66,71,67,69,71,74,78,67,68,67,65,71,70,75,83,64,65,68,65,69,73,72,77,58,65,62,71,66,68,72,71,61,69,65,65,68,68,73,71);
		wait for 10 ns;
		t_blur_matrix_int <= (81,82,83,85,83,87,82,85,78,83,80,83,84,85,87,83,79,84,83,83,84,83,81,134,83,82,82,85,86,83,89,189,80,80,83,87,91,90,98,163,81,82,82,84,96,109,104,108,73,79,78,101,123,127,111,110,75,76,84,120,128,128,121,117);
		wait for 10 ns;
		t_blur_matrix_int <= (81,91,118,56,86,132,143,76,90,91,149,91,89,105,156,102,174,132,96,15,20,23,39,89,136,60,32,11,13,12,38,120,134,54,28,21,11,16,76,129,133,87,31,19,12,17,76,110,123,86,30,60,47,16,79,98,133,158,110,123,108,70,98,85);
		wait for 10 ns;
		t_blur_matrix_int <= (86,94,96,109,92,84,91,70,86,94,104,96,84,92,86,34,106,100,99,85,76,80,58,22,159,167,85,66,68,51,19,30,148,139,82,43,45,43,28,41,91,57,68,32,56,41,29,61,97,50,53,55,33,26,45,77,106,61,40,33,24,36,55,96);
		wait for 10 ns;
		t_blur_matrix_int <= (30,28,83,32,10,12,87,56,20,44,89,16,10,17,89,74,46,58,74,9,13,33,99,56,63,79,36,16,16,55,114,46,66,93,17,15,34,67,113,53,65,31,17,24,65,59,74,71,54,22,25,63,77,22,52,103,48,39,47,88,49,8,22,90);
		wait for 10 ns;
		t_blur_matrix_int <= (29,17,26,20,40,35,77,60,15,14,17,16,43,69,59,49,10,18,26,34,38,28,27,29,8,24,16,21,25,26,30,33,8,16,13,34,50,41,25,46,9,15,29,56,37,33,54,45,18,17,21,40,29,15,20,49,37,19,23,61,21,16,12,40);
		wait for 10 ns;
		t_blur_matrix_int <= (42,25,11,18,31,13,25,64,33,16,19,17,29,20,40,49,16,13,18,18,25,24,39,24,19,20,30,21,21,36,45,34,32,20,28,18,17,15,44,71,49,21,25,13,15,10,17,55,75,34,12,11,14,16,13,34,81,45,16,10,14,22,14,15);
		wait for 10 ns;
		t_blur_matrix_int <= (13,27,74,30,19,61,47,16,10,20,85,21,17,71,18,30,10,46,79,18,37,54,37,17,23,46,60,29,48,23,10,11,24,60,40,37,40,13,13,43,62,81,16,56,24,8,18,97,55,88,21,42,8,6,62,132,15,32,51,9,8,34,124,91);
		wait for 10 ns;
		t_blur_matrix_int <= (18,11,51,112,75,69,128,161,20,27,113,96,59,120,170,143,18,92,124,68,93,175,153,146,68,123,76,79,155,160,150,161,121,96,72,139,156,153,162,169,127,76,127,174,145,156,167,183,99,106,171,151,151,164,176,190,89,167,159,150,160,177,186,189);
		wait for 10 ns;
		t_blur_matrix_int <= (140,143,146,137,140,156,178,180,152,160,153,140,137,157,177,178,162,169,152,132,129,155,179,182,172,180,141,132,137,167,180,186,185,172,135,132,150,174,178,186,188,154,129,144,165,181,188,178,179,140,133,159,180,189,172,94,166,147,150,173,192,158,74,65);
		wait for 10 ns;
		t_blur_matrix_int <= (171,175,167,161,169,159,146,131,176,178,170,170,162,124,84,97,186,178,180,159,79,42,58,74,185,184,143,72,67,74,76,69,182,130,91,101,115,113,114,104,113,83,101,113,123,116,112,130,81,92,92,107,105,106,72,119,74,70,72,79,79,75,26,67);
		wait for 10 ns;
		t_blur_matrix_int <= (125,134,137,139,138,138,141,142,113,120,126,134,139,141,145,149,80,94,103,105,115,126,141,147,63,66,53,62,75,86,109,130,93,81,60,33,35,36,51,70,127,107,88,74,53,46,35,32,130,116,90,95,63,61,55,49,115,80,61,65,68,88,68,75);
		wait for 10 ns;
		t_blur_matrix_int <= (148,156,153,152,156,155,152,158,153,153,155,158,156,154,155,161,150,155,159,157,152,153,152,153,144,154,161,156,154,151,154,148,105,129,151,151,153,158,152,150,40,67,112,139,145,145,139,146,46,52,69,104,137,138,139,140,65,68,67,90,116,124,128,137);
		wait for 10 ns;
		t_blur_matrix_int <= (168,171,177,183,181,180,179,184,163,168,174,179,180,179,180,179,161,161,170,180,182,179,175,173,154,163,169,176,178,178,170,171,151,155,168,175,177,179,167,172,151,155,167,172,173,173,170,169,143,149,163,167,176,176,170,169,136,145,163,172,177,179,175,170);
		wait for 10 ns;
		t_blur_matrix_int <= (186,187,188,192,193,196,197,200,181,185,188,189,189,192,195,200,180,180,185,187,186,190,194,194,176,178,182,186,186,189,193,191,173,175,177,187,184,185,184,172,180,177,171,177,165,150,118,85,173,167,162,162,123,83,54,60,174,164,147,126,89,87,79,85);
		wait for 10 ns;
		t_blur_matrix_int <= (198,198,193,169,122,74,55,36,197,192,192,171,130,78,43,27,194,189,178,154,118,67,30,20,186,174,145,117,82,51,28,20,143,113,87,74,60,40,28,23,68,52,50,57,70,67,62,49,73,74,85,86,100,75,68,52,82,56,56,72,64,48,46,39);
		wait for 10 ns;
		t_blur_matrix_int <= (17,13,17,19,42,46,123,158,16,12,16,15,28,34,121,163,20,11,12,15,28,38,102,165,14,11,13,12,31,46,74,170,12,12,16,19,28,34,62,165,20,18,18,16,22,37,58,165,30,26,15,16,18,38,47,157,32,39,19,19,22,44,44,153);
		wait for 10 ns;
		t_blur_matrix_int <= (100,44,37,25,35,41,33,37,112,43,43,29,43,42,31,31,124,49,33,32,37,35,40,36,128,75,29,25,45,36,33,31,137,89,27,23,34,39,42,34,131,102,37,29,29,49,44,39,135,96,45,23,28,50,31,34,137,94,64,20,23,47,32,40);
		wait for 10 ns;
		t_blur_matrix_int <= (33,38,40,36,28,27,28,26,36,36,40,31,25,21,29,25,41,48,49,33,23,21,26,24,39,45,37,26,20,23,21,29,39,34,30,31,28,23,25,24,43,35,29,20,27,23,22,23,40,40,28,24,28,24,27,27,40,34,23,22,22,25,27,29);
		wait for 10 ns;
		t_blur_matrix_int <= (23,28,22,22,20,43,90,116,27,32,24,18,31,65,98,114,25,30,22,24,33,78,109,117,27,26,19,23,46,87,112,118,34,24,24,23,57,99,115,112,32,29,26,27,69,112,115,108,30,30,29,36,82,113,116,107,27,21,32,51,98,114,113,103);
		wait for 10 ns;
		t_blur_matrix_int <= (116,109,104,123,136,145,143,145,114,107,111,128,139,143,145,143,110,104,114,133,141,143,141,138,111,102,121,138,144,141,141,141,106,108,128,140,146,143,137,140,104,116,131,142,141,142,139,139,105,124,138,142,143,139,138,141,106,128,139,140,137,137,135,134);
		wait for 10 ns;
		t_blur_matrix_int <= (145,144,141,143,143,146,142,147,145,143,143,142,140,144,145,144,141,142,139,141,143,142,138,143,138,138,140,139,139,139,140,139,138,139,137,139,136,138,136,136,138,137,138,138,138,138,136,135,137,136,136,138,136,135,134,137,137,134,135,134,137,135,134,135);
		wait for 10 ns;
		t_blur_matrix_int <= (148,150,147,149,148,141,140,139,147,146,151,148,144,145,141,138,143,145,145,145,146,144,138,137,138,141,144,143,141,144,144,136,137,139,138,140,141,142,141,136,135,138,139,140,140,141,140,135,135,134,137,137,138,141,137,136,135,137,137,139,140,139,138,136);
		wait for 10 ns;
		t_blur_matrix_int <= (136,131,130,131,128,130,125,124,138,141,135,133,131,132,127,127,138,138,136,139,134,133,133,132,133,134,140,137,139,137,137,134,134,135,135,138,135,135,134,138,138,136,134,136,137,136,139,135,135,136,133,134,136,135,138,140,136,135,134,134,134,134,131,136);
		wait for 10 ns;
		t_blur_matrix_int <= (125,121,124,122,123,123,120,122,125,125,125,123,121,121,123,122,129,128,127,128,128,126,124,121,132,130,134,127,129,127,122,123,135,138,133,135,131,130,125,124,136,137,138,137,135,132,129,129,136,137,138,134,134,133,132,133,138,139,139,137,139,134,129,131);
		wait for 10 ns;
		t_blur_matrix_int <= (122,124,126,127,126,126,128,132,118,121,122,120,119,124,123,125,122,123,122,121,120,117,117,117,120,120,120,119,118,119,114,113,123,122,125,119,119,113,111,111,123,125,123,119,117,114,115,110,131,127,126,120,117,113,113,110,134,134,127,123,118,117,117,110);
		wait for 10 ns;
		t_blur_matrix_int <= (64,69,69,71,70,68,66,65,64,72,68,68,65,67,64,67,62,68,67,62,68,64,60,60,62,60,65,60,60,64,58,59,62,69,66,61,59,62,59,57,67,65,65,62,63,64,60,59,65,65,71,60,68,61,64,60,70,66,65,64,65,64,66,56);
		wait for 10 ns;
		t_blur_matrix_int <= (67,60,60,50,49,63,87,100,61,65,56,55,49,63,86,102,60,60,53,48,47,56,80,100,57,57,52,44,42,53,80,97,58,52,48,47,40,52,77,101,55,51,49,44,39,56,80,102,56,58,50,44,37,52,78,97,61,56,48,42,38,51,76,97);
		wait for 10 ns;
		t_blur_matrix_int <= (117,128,139,150,156,155,152,155,117,125,140,147,152,157,155,159,116,128,142,145,153,155,157,158,115,125,141,153,154,155,154,158,114,129,142,153,156,152,156,155,114,130,142,155,157,157,153,158,114,129,141,151,156,156,158,160,114,128,140,151,158,157,156,162);
		wait for 10 ns;
		t_blur_matrix_int <= (156,156,154,142,135,124,110,81,156,154,152,146,134,120,102,82,156,154,153,141,131,119,109,82,155,156,154,143,132,120,101,82,155,158,152,145,132,118,102,83,160,159,157,153,132,119,100,82,163,161,156,146,134,117,102,83,162,159,156,151,136,117,100,83);
		wait for 10 ns;
		t_blur_matrix_int <= (60,43,40,48,51,51,64,63,59,51,42,42,49,52,57,59,59,46,37,45,50,54,54,53,56,40,39,39,50,54,57,57,57,42,40,44,50,53,59,62,57,40,41,48,51,57,66,60,61,43,42,48,49,61,64,64,63,49,43,51,54,58,64,65);
		wait for 10 ns;
		t_blur_matrix_int <= (65,66,66,69,65,63,65,65,63,69,66,67,65,65,65,60,64,60,72,67,63,62,61,64,61,61,62,64,61,60,62,58,65,62,62,62,61,66,60,65,63,65,65,63,61,66,68,66,68,67,66,69,68,70,70,64,68,70,67,69,73,63,70,73);
		wait for 10 ns;
		t_blur_matrix_int <= (64,64,57,62,66,64,69,77,62,62,66,60,58,60,82,123,62,62,60,53,52,70,129,153,61,57,56,46,47,132,184,180,58,55,53,51,48,143,170,185,63,57,56,50,33,90,162,165,69,62,61,39,15,76,149,50,89,49,31,29,20,28,141,98);
		wait for 10 ns;
		t_blur_matrix_int <= (89,110,112,115,127,130,127,123,140,139,113,119,122,127,124,123,198,122,107,118,119,123,125,123,186,89,111,113,118,127,127,97,128,94,108,115,124,126,113,67,168,131,117,117,119,120,107,91,95,175,173,137,127,122,80,44,151,169,200,209,173,84,24,18);
		wait for 10 ns;
		t_blur_matrix_int <= (126,150,137,142,137,87,46,35,127,121,77,84,109,60,16,14,122,101,67,28,59,45,12,9,112,94,45,43,28,15,10,13,105,92,43,36,14,20,21,61,123,58,23,22,15,31,70,67,47,21,12,16,23,72,72,29,18,16,12,23,60,58,31,34);
		wait for 10 ns;
		t_blur_matrix_int <= (32,22,50,34,40,58,93,61,8,24,55,55,59,81,106,39,20,71,88,51,57,98,49,66,85,95,38,25,89,42,26,61,87,34,16,73,56,12,15,53,19,18,50,48,33,17,20,57,16,51,44,28,55,20,28,69,28,46,43,33,46,42,48,91);
		wait for 10 ns;
		t_blur_matrix_int <= (28,54,51,91,38,8,17,59,35,71,52,96,35,16,24,52,48,63,66,110,34,17,21,50,65,53,93,109,27,11,29,48,95,69,88,67,24,16,27,30,100,59,91,61,27,21,21,17,94,58,117,62,21,20,22,21,98,60,123,71,19,19,25,22);
		wait for 10 ns;
		t_blur_matrix_int <= (57,17,26,65,18,14,12,27,49,24,22,76,19,12,11,17,16,45,26,87,20,16,12,10,19,37,39,94,33,22,20,15,15,23,16,79,61,21,19,18,16,19,15,49,87,34,19,10,23,16,13,32,99,40,18,19,34,18,18,22,65,28,20,25);
		wait for 10 ns;
		t_blur_matrix_int <= (65,80,21,19,19,16,18,20,30,95,76,28,17,18,19,21,11,44,94,90,42,10,12,18,15,18,52,85,72,56,27,13,18,20,24,28,19,40,54,24,15,17,28,22,14,28,28,14,16,18,30,16,12,16,12,15,18,16,26,20,15,10,15,23);
		wait for 10 ns;
		t_blur_matrix_int <= (16,13,22,19,9,89,119,74,13,13,16,6,50,135,89,108,17,15,10,18,110,110,87,169,10,10,9,71,131,71,139,178,9,8,24,120,91,93,179,152,29,39,78,118,68,162,172,150,12,40,92,62,108,163,135,128,26,89,85,72,152,138,146,160);
		wait for 10 ns;
		t_blur_matrix_int <= (144,169,150,155,169,186,192,186,180,152,157,163,178,191,189,178,160,148,161,167,180,193,185,178,149,156,161,169,188,193,187,179,154,165,164,173,197,190,185,192,163,171,175,190,194,192,191,171,145,165,186,192,191,188,177,90,175,186,191,188,188,178,92,78);
		wait for 10 ns;
		t_blur_matrix_int <= (170,156,168,189,145,54,53,54,173,169,188,132,42,42,38,31,179,182,140,42,31,29,19,20,187,144,42,40,33,23,17,20,154,55,52,43,25,17,11,26,70,64,53,32,21,19,14,35,71,82,73,56,49,26,14,38,84,94,92,89,81,59,16,25);
		wait for 10 ns;
		t_blur_matrix_int <= (50,59,36,33,35,30,16,29,22,26,22,23,18,18,20,24,21,22,24,18,15,16,16,38,19,20,18,17,15,23,28,70,48,29,35,28,9,31,47,56,73,48,46,61,26,40,68,39,72,87,40,54,58,55,31,97,68,87,81,46,31,42,94,176);
		wait for 10 ns;
		t_blur_matrix_int <= (46,24,19,26,52,86,64,92,26,24,15,10,14,27,85,106,67,57,27,17,14,12,27,74,150,150,89,35,13,12,13,41,173,189,167,127,43,25,58,41,174,189,189,177,109,36,76,63,198,199,198,192,147,64,53,82,193,193,189,177,135,94,65,86);
		wait for 10 ns;
		t_blur_matrix_int <= (85,82,80,90,100,116,127,129,92,90,88,92,104,110,118,126,101,96,90,91,99,106,114,118,89,97,90,89,98,101,109,118,79,88,80,86,95,101,111,110,63,81,75,84,90,98,103,107,57,71,74,80,84,94,99,112,75,74,86,78,84,94,103,112);
		wait for 10 ns;
		t_blur_matrix_int <= (127,142,159,174,176,181,177,174,130,140,160,174,177,182,185,182,128,140,162,175,187,187,191,186,125,137,161,177,193,194,198,174,125,137,156,185,199,204,194,111,122,144,165,190,207,208,152,62,129,145,171,194,206,197,111,61,130,146,181,204,209,187,83,76);
		wait for 10 ns;
		t_blur_matrix_int <= (172,166,134,109,96,87,51,41,174,150,107,60,38,27,19,22,159,91,40,28,25,29,22,39,80,22,24,18,28,34,50,86,31,23,22,19,25,41,119,91,39,30,48,24,26,44,62,83,81,38,69,61,53,64,36,115,107,87,51,65,65,46,89,159);
		wait for 10 ns;
		t_blur_matrix_int <= (25,20,22,30,31,34,38,32,21,17,18,23,29,26,28,34,39,24,20,21,31,32,26,27,106,63,20,13,19,25,26,25,143,101,41,18,13,26,23,26,155,123,57,28,18,25,18,22,149,121,65,31,15,15,11,18,148,113,59,29,19,15,17,18);
		wait for 10 ns;
		t_blur_matrix_int <= (43,20,18,11,21,48,37,151,33,13,18,12,14,50,30,147,19,19,17,14,22,42,28,137,15,21,20,13,20,46,23,133,19,19,19,11,26,45,18,129,20,18,30,21,23,51,18,132,18,17,17,16,29,51,17,124,16,16,15,15,41,48,22,117);
		wait for 10 ns;
		t_blur_matrix_int <= (144,87,70,27,22,50,33,39,153,93,68,47,21,43,41,35,152,92,71,43,35,42,38,36,161,94,65,38,32,46,45,34,157,92,66,56,40,51,38,36,156,111,51,68,42,59,34,34,161,121,50,70,46,64,30,34,160,123,49,64,53,59,31,29);
		wait for 10 ns;
		t_blur_matrix_int <= (33,27,24,22,21,24,23,27,37,27,19,22,25,23,26,29,30,21,21,24,23,24,26,32,28,20,18,23,22,24,30,24,30,18,20,21,31,30,22,20,26,20,27,24,22,25,19,20,22,21,24,27,28,27,22,26,23,28,26,24,36,24,19,19);
		wait for 10 ns;
		t_blur_matrix_int <= (23,15,29,72,112,119,112,103,25,12,27,84,116,115,109,106,23,16,35,93,121,112,110,115,23,23,58,107,120,118,111,122,20,33,80,114,122,115,112,128,30,47,94,118,116,115,115,131,24,63,106,119,116,110,120,133,25,77,114,121,117,115,127,137);
		wait for 10 ns;
		t_blur_matrix_int <= (117,133,141,141,138,138,137,133,121,136,138,139,138,138,136,134,132,142,139,139,136,135,134,130,138,141,136,139,137,133,135,132,138,140,137,135,137,136,135,129,141,137,137,135,136,136,133,132,139,136,138,137,135,137,132,132,140,138,135,134,132,136,130,133);
		wait for 10 ns;
		t_blur_matrix_int <= (134,134,138,137,135,134,132,131,136,133,130,136,136,135,133,136,135,132,131,132,134,130,135,136,131,130,130,134,130,131,131,137,136,132,132,131,130,132,132,133,130,131,129,132,134,131,127,131,132,132,131,131,126,129,131,132,128,132,130,131,133,131,128,131);
		wait for 10 ns;
		t_blur_matrix_int <= (135,136,136,138,136,137,137,134,135,135,137,136,138,138,139,132,132,131,133,135,134,135,135,132,131,131,135,137,135,131,135,132,131,131,133,130,130,133,134,134,130,131,131,129,129,132,127,133,131,133,130,131,137,131,132,130,128,133,133,129,129,130,132,130);
		wait for 10 ns;
		t_blur_matrix_int <= (133,133,131,134,135,138,134,136,133,134,136,131,134,133,133,134,135,133,133,135,132,135,131,130,133,132,136,134,131,131,134,130,134,132,131,135,131,131,129,128,132,132,131,130,127,129,126,127,131,128,127,127,129,130,125,126,129,132,128,124,128,128,125,129);
		wait for 10 ns;
		t_blur_matrix_int <= (137,136,138,136,134,130,128,126,134,135,134,136,132,132,127,128,134,132,134,132,128,126,127,124,131,132,132,128,126,124,124,121,130,133,130,125,124,121,120,118,128,127,125,124,122,121,122,118,125,125,121,124,117,120,117,111,123,127,120,115,116,117,113,109);
		wait for 10 ns;
		t_blur_matrix_int <= (129,128,125,126,121,118,119,114,124,127,125,123,122,119,116,115,125,122,122,120,120,119,119,114,121,116,117,118,119,116,116,113,116,118,112,117,115,113,114,111,115,110,113,111,110,107,109,117,109,110,105,109,111,121,129,140,110,107,114,121,130,138,147,158);
		wait for 10 ns;
		t_blur_matrix_int <= (64,69,68,64,65,65,65,57,68,69,69,66,64,66,63,56,73,72,68,67,74,69,61,56,67,67,72,72,66,68,59,56,68,70,70,67,66,67,59,55,66,72,66,67,63,61,56,53,68,66,63,59,61,57,54,50,68,60,57,56,60,53,49,45);
		wait for 10 ns;
		t_blur_matrix_int <= (60,57,49,42,35,54,76,96,56,57,54,40,37,51,78,100,56,49,46,45,36,49,77,97,51,51,46,38,35,47,71,97,49,54,46,41,37,43,73,97,50,52,47,37,29,45,69,94,49,47,41,29,22,37,67,96,49,46,38,30,29,35,64,95);
		wait for 10 ns;
		t_blur_matrix_int <= (116,126,141,149,158,158,161,159,115,128,138,150,155,158,161,159,114,129,143,149,153,157,160,161,115,130,140,152,155,157,161,166,113,127,142,149,155,160,159,163,113,128,141,149,157,157,162,161,113,126,138,146,153,160,162,161,113,124,140,149,155,158,162,162);
		wait for 10 ns;
		t_blur_matrix_int <= (159,158,158,150,135,120,100,81,165,158,160,150,137,122,102,86,161,163,160,153,139,123,105,85,168,163,165,151,143,125,103,87,162,163,163,153,143,124,106,87,163,163,158,156,140,126,108,90,163,163,163,154,139,126,109,89,163,162,163,155,141,126,106,89);
		wait for 10 ns;
		t_blur_matrix_int <= (62,47,50,51,57,62,66,70,64,51,53,53,55,60,64,69,63,49,48,55,60,62,69,71,66,46,48,54,62,67,68,68,68,45,45,49,57,62,65,70,65,44,43,53,59,61,68,69,62,46,46,54,56,60,64,69,64,51,41,50,56,60,63,72);
		wait for 10 ns;
		t_blur_matrix_int <= (70,74,71,72,71,69,63,51,71,75,72,72,77,92,23,16,77,76,79,75,93,88,14,13,76,74,75,70,87,104,24,43,75,81,73,71,73,121,97,111,72,70,71,70,68,95,127,119,72,74,71,70,73,77,107,138,76,76,75,74,74,86,92,94);
		wait for 10 ns;
		t_blur_matrix_int <= (40,23,48,35,60,94,152,129,16,29,82,107,126,126,147,170,43,74,133,130,119,121,113,136,98,108,141,110,105,106,99,126,114,99,116,137,93,56,43,52,143,141,111,82,51,50,43,56,121,89,87,73,39,33,58,74,79,81,69,46,62,76,79,49);
		wait for 10 ns;
		t_blur_matrix_int <= (148,184,238,221,113,32,48,15,158,201,147,60,26,28,72,24,165,105,32,31,20,22,71,79,82,38,45,32,24,23,30,102,70,50,27,15,19,20,17,52,64,38,19,14,36,22,23,27,45,31,13,23,56,28,44,50,25,27,20,29,65,43,74,91);
		wait for 10 ns;
		t_blur_matrix_int <= (17,14,18,52,74,59,53,39,23,40,79,111,91,64,15,14,78,87,69,47,70,31,11,15,94,43,29,85,73,19,18,21,122,107,88,114,75,75,34,31,54,124,118,104,104,82,33,25,71,78,70,68,78,48,19,13,98,62,28,53,81,34,14,17);
		wait for 10 ns;
		t_blur_matrix_int <= (20,47,54,60,58,67,48,98,12,65,26,66,54,49,55,107,27,87,24,71,53,44,55,88,25,82,36,65,75,23,49,88,13,67,38,49,88,43,54,78,16,43,54,37,79,83,69,50,15,32,50,39,33,89,97,79,26,32,64,64,30,33,113,133);
		wait for 10 ns;
		t_blur_matrix_int <= (85,48,115,88,29,30,20,18,103,40,131,99,61,35,35,18,118,70,135,81,65,49,57,19,93,90,115,68,85,114,25,13,80,108,109,107,123,41,13,27,50,89,86,122,82,61,45,34,86,71,68,85,48,77,30,24,96,45,64,65,140,56,18,21);
		wait for 10 ns;
		t_blur_matrix_int <= (29,19,14,18,35,23,28,28,19,10,14,21,23,21,31,25,19,13,19,20,21,19,20,17,18,22,23,16,20,20,17,18,23,19,25,23,17,24,20,21,14,20,21,20,19,20,25,22,20,17,20,17,18,16,25,23,23,20,25,17,17,18,22,28);
		wait for 10 ns;
		t_blur_matrix_int <= (18,17,22,18,14,12,8,26,21,23,35,18,16,11,12,30,22,27,22,12,10,9,10,77,27,25,14,12,8,10,41,120,28,23,16,9,6,16,103,112,18,19,14,13,8,57,126,82,23,25,17,12,26,111,101,69,26,29,23,21,69,122,68,87);
		wait for 10 ns;
		t_blur_matrix_int <= (67,118,66,129,167,130,158,168,114,77,93,184,154,148,165,176,114,61,149,172,147,157,173,186,73,89,173,144,155,168,178,189,71,128,153,148,164,167,186,195,92,168,148,157,171,183,196,192,125,162,163,170,180,195,196,104,156,159,172,178,190,202,127,33);
		wait for 10 ns;
		t_blur_matrix_int <= (183,188,191,187,170,89,80,86,192,193,190,170,79,75,87,90,194,191,173,75,67,80,95,93,194,176,74,59,73,91,98,100,181,78,48,65,79,92,98,103,83,48,58,73,84,90,102,111,37,56,72,75,83,98,97,107,46,63,75,81,86,93,103,105);
		wait for 10 ns;
		t_blur_matrix_int <= (82,87,104,105,100,83,54,50,95,90,106,113,110,104,93,72,100,98,105,109,109,113,107,91,109,102,110,111,112,110,112,113,113,111,115,115,120,113,107,111,117,122,121,119,122,123,123,121,117,121,124,124,131,133,132,132,117,119,126,127,134,142,134,138);
		wait for 10 ns;
		t_blur_matrix_int <= (63,81,101,96,90,117,166,183,66,68,83,99,115,126,140,155,98,91,72,81,62,91,104,102,113,98,84,91,68,96,104,99,119,107,106,103,95,99,107,107,116,109,113,111,108,111,112,123,128,120,123,129,122,131,135,138,148,149,140,138,140,138,149,151);
		wait for 10 ns;
		t_blur_matrix_int <= (190,196,192,158,108,115,91,78,164,164,159,157,133,111,96,93,109,99,125,145,150,156,140,109,89,92,122,120,130,131,117,102,104,119,126,128,124,116,121,118,123,130,136,138,131,135,136,111,142,144,139,143,134,141,132,108,147,145,139,146,138,140,124,105);
		wait for 10 ns;
		t_blur_matrix_int <= (95,80,78,84,90,91,96,105,95,87,81,80,90,93,87,111,86,86,85,90,88,92,93,106,85,83,92,95,88,90,87,106,88,86,97,98,92,90,86,95,95,95,99,99,92,87,88,90,94,99,107,99,87,90,89,89,101,111,106,99,91,91,90,89);
		wait for 10 ns;
		t_blur_matrix_int <= (126,152,189,212,210,173,79,60,126,153,185,213,210,169,106,78,121,152,182,213,213,176,150,142,119,141,176,210,216,181,145,127,120,138,177,207,217,190,154,136,115,141,175,201,214,194,169,154,113,137,167,201,216,196,175,163,111,141,168,200,213,202,176,165);
		wait for 10 ns;
		t_blur_matrix_int <= (91,112,95,72,77,108,161,161,75,88,115,115,122,137,145,133,128,112,118,99,94,108,113,73,115,107,104,85,82,85,80,57,125,109,101,94,98,92,94,79,137,127,114,106,104,94,89,86,142,131,127,120,112,94,93,94,152,137,129,124,119,105,99,94);
		wait for 10 ns;
		t_blur_matrix_int <= (146,103,56,27,24,21,16,23,112,71,42,15,35,33,24,26,52,36,28,28,55,46,24,25,41,39,53,52,51,40,21,23,62,53,63,63,62,48,21,25,72,69,71,73,65,49,26,31,86,79,81,79,73,57,29,29,88,82,82,75,71,59,27,27);
		wait for 10 ns;
		t_blur_matrix_int <= (25,17,30,21,45,42,25,99,23,24,34,27,48,43,25,99,25,19,34,25,48,35,21,92,17,13,25,31,54,40,24,86,13,16,19,25,45,39,19,87,13,19,22,31,42,36,23,82,15,20,23,34,43,38,20,78,19,22,26,35,37,30,17,70);
		wait for 10 ns;
		t_blur_matrix_int <= (163,131,55,62,61,59,38,21,157,144,70,60,72,36,33,28,149,146,86,51,66,44,36,20,148,157,99,45,72,41,28,22,142,164,109,49,63,37,23,24,141,160,111,49,50,35,23,29,141,166,120,54,53,40,25,26,142,164,130,50,48,33,18,31);
		wait for 10 ns;
		t_blur_matrix_int <= (24,24,20,21,29,27,24,18,17,22,17,22,29,29,17,27,24,24,22,22,34,27,24,59,25,26,16,29,29,23,24,56,21,17,18,40,27,19,21,61,27,22,25,39,23,16,23,73,21,14,24,28,21,18,32,87,20,16,26,27,17,16,43,95);
		wait for 10 ns;
		t_blur_matrix_int <= (40,90,116,116,112,116,131,141,54,102,120,114,110,122,136,140,75,105,116,108,111,124,138,138,92,116,113,108,118,132,141,140,107,113,109,105,120,138,141,137,112,111,110,107,125,137,136,136,115,114,109,113,127,137,138,133,113,108,111,118,136,139,134,135);
		wait for 10 ns;
		t_blur_matrix_int <= (137,137,135,135,134,132,132,131,135,133,137,134,131,134,131,131,134,136,135,134,129,131,130,127,137,134,132,132,132,132,132,131,136,132,134,131,132,128,132,128,135,130,133,133,131,127,126,131,136,136,129,131,129,130,129,131,136,132,131,130,130,129,128,131);
		wait for 10 ns;
		t_blur_matrix_int <= (130,130,129,133,143,133,131,133,126,131,131,133,140,147,131,133,128,130,129,134,140,145,130,131,132,129,127,130,130,129,130,134,133,131,132,132,128,129,130,129,133,130,129,129,128,128,129,129,131,130,128,131,133,128,128,129,127,134,132,132,129,126,128,130);
		wait for 10 ns;
		t_blur_matrix_int <= (131,133,135,135,133,131,131,129,129,132,134,133,129,130,128,127,130,132,133,135,135,130,128,125,128,127,130,133,129,130,129,125,131,129,129,130,131,127,126,126,129,131,130,132,125,123,125,122,129,127,129,129,126,124,124,123,127,126,125,128,126,124,124,120);
		wait for 10 ns;
		t_blur_matrix_int <= (129,130,128,127,128,123,124,120,127,125,125,124,121,124,121,120,125,124,124,118,116,120,120,115,123,124,120,121,119,117,113,114,122,126,120,117,119,117,113,116,121,118,121,122,117,113,115,108,120,121,119,121,113,110,109,114,123,122,119,115,112,111,114,140);
		wait for 10 ns;
		t_blur_matrix_int <= (121,121,119,121,112,113,110,107,116,118,120,115,114,109,116,124,112,117,116,116,113,123,134,147,115,112,115,121,134,145,157,165,111,113,126,141,155,164,173,177,116,130,151,165,172,178,183,181,136,155,171,181,183,184,184,184,159,171,181,187,187,186,185,181);
		wait for 10 ns;
		t_blur_matrix_int <= (116,126,133,143,150,157,162,171,141,147,152,163,166,170,173,178,159,164,168,171,176,174,176,180,170,173,179,178,180,176,175,176,180,179,179,180,179,180,176,177,180,182,178,178,179,179,177,178,182,182,181,178,178,178,180,178,180,181,179,178,179,179,177,179);
		wait for 10 ns;
		t_blur_matrix_int <= (60,59,58,57,52,53,52,46,58,60,69,58,56,52,53,52,56,58,65,55,52,48,47,47,54,52,59,53,47,44,53,45,52,49,47,49,46,40,46,48,50,48,48,46,46,43,43,41,50,48,44,42,40,42,38,39,45,44,46,43,47,46,45,39);
		wait for 10 ns;
		t_blur_matrix_int <= (46,46,34,29,27,42,64,93,45,44,35,28,27,40,62,90,43,40,35,29,22,40,72,91,42,38,38,28,24,39,67,92,41,41,33,27,29,32,64,93,43,41,34,32,26,35,63,91,38,36,31,28,22,36,58,92,36,37,31,22,24,33,58,91);
		wait for 10 ns;
		t_blur_matrix_int <= (108,124,138,147,154,159,158,159,109,129,141,149,157,157,158,160,112,127,137,148,154,157,160,160,115,125,141,148,155,155,159,156,111,125,143,150,154,156,158,159,108,123,140,146,153,154,161,160,112,124,136,147,150,156,158,155,114,124,134,145,147,153,154,151);
		wait for 10 ns;
		t_blur_matrix_int <= (165,161,162,153,140,126,110,89,163,160,160,151,140,127,108,84,161,161,160,153,137,125,107,89,160,166,162,150,139,128,109,87,164,159,159,152,139,121,108,83,158,159,156,150,137,120,107,90,154,155,152,149,136,125,108,91,156,156,156,149,139,124,107,90);
		wait for 10 ns;
		t_blur_matrix_int <= (67,48,45,49,57,60,64,66,62,48,44,50,59,58,62,62,65,42,42,49,54,55,62,68,60,48,43,48,54,57,68,97,67,47,41,53,52,59,71,78,64,48,45,52,56,65,63,75,64,44,45,49,57,56,68,70,62,42,44,50,61,71,63,67);
		wait for 10 ns;
		t_blur_matrix_int <= (72,76,74,78,77,86,80,76,67,72,81,92,109,120,126,137,78,105,132,122,127,112,112,116,105,91,81,86,101,95,100,74,71,76,78,86,100,78,70,61,75,76,78,82,95,61,58,52,70,70,77,78,79,42,61,100,70,73,73,75,78,74,134,121);
		wait for 10 ns;
		t_blur_matrix_int <= (109,119,100,118,137,117,74,35,137,146,120,95,85,63,41,33,112,59,32,39,61,41,31,37,55,34,41,58,55,35,38,32,71,63,63,63,47,41,28,32,53,73,77,49,77,49,26,44,109,96,47,60,80,52,53,88,88,49,59,85,72,44,93,78);
		wait for 10 ns;
		t_blur_matrix_int <= (31,30,26,41,83,50,100,87,37,44,32,60,77,53,95,87,38,36,38,71,65,59,94,63,39,41,63,60,55,90,88,117,45,72,87,32,53,108,118,98,78,93,42,30,67,126,80,85,80,40,24,30,45,106,97,75,37,37,39,37,28,66,118,66);
		wait for 10 ns;
		t_blur_matrix_int <= (83,55,53,103,63,14,15,17,65,88,98,70,24,14,15,14,101,109,73,41,23,25,20,16,108,101,31,23,29,21,20,24,41,47,49,24,28,19,22,21,42,56,49,27,19,19,22,30,62,39,39,24,20,23,29,28,84,28,38,31,26,25,35,21);
		wait for 10 ns;
		t_blur_matrix_int <= (20,38,74,100,63,49,51,67,25,25,31,66,78,88,92,76,16,18,23,43,50,56,95,107,23,20,23,27,46,63,31,44,19,19,31,23,22,46,58,31,26,23,28,24,25,36,30,27,28,24,26,24,28,32,29,20,23,23,20,18,19,35,80,19);
		wait for 10 ns;
		t_blur_matrix_int <= (100,70,97,140,102,35,37,33,61,125,139,92,46,92,72,57,106,53,25,19,50,117,103,80,67,19,13,20,59,110,110,79,53,20,10,16,69,100,113,81,56,19,7,18,67,98,100,127,45,23,10,32,68,94,74,137,15,32,18,15,66,89,62,80);
		wait for 10 ns;
		t_blur_matrix_int <= (25,20,26,25,21,17,23,25,51,15,23,26,17,21,21,21,51,25,24,21,25,24,22,22,43,24,18,22,23,19,21,20,74,25,22,19,21,14,23,18,82,25,15,15,14,12,18,11,118,56,12,16,12,10,11,7,151,120,50,18,12,15,11,13);
		wait for 10 ns;
		t_blur_matrix_int <= (26,22,24,30,120,95,74,138,20,17,18,82,123,69,87,165,23,20,31,125,98,78,124,167,15,21,77,122,83,92,157,161,12,37,126,101,84,129,178,176,8,77,115,80,92,176,175,181,28,120,95,83,119,178,180,188,68,114,73,90,163,177,189,203);
		wait for 10 ns;
		t_blur_matrix_int <= (159,169,178,184,193,155,29,38,158,178,181,196,180,45,23,38,174,183,192,199,72,13,26,45,180,186,204,121,14,15,28,57,176,191,161,23,16,22,34,56,179,191,56,17,22,21,38,59,199,111,23,21,27,25,34,57,170,29,12,24,29,22,35,55);
		wait for 10 ns;
		t_blur_matrix_int <= (52,69,76,85,87,90,105,102,57,75,78,82,89,91,97,104,61,75,79,85,87,90,99,106,67,80,84,86,89,93,94,102,72,82,81,86,87,86,96,104,74,79,82,88,90,91,94,94,71,83,81,83,91,96,94,95,68,78,84,87,88,93,93,102);
		wait for 10 ns;
		t_blur_matrix_int <= (112,120,125,127,133,145,135,140,112,120,120,127,132,142,145,143,112,118,118,126,132,139,148,147,111,111,120,124,131,139,141,148,107,115,120,122,126,135,145,150,102,111,114,114,124,132,140,143,104,110,110,114,122,123,129,136,103,110,114,116,120,122,127,135);
		wait for 10 ns;
		t_blur_matrix_int <= (148,152,147,143,142,143,148,148,149,152,147,157,151,152,147,143,149,158,152,144,156,154,157,155,151,156,156,153,154,154,152,154,152,157,155,156,161,156,153,148,149,150,156,155,161,162,150,147,139,147,154,154,153,161,151,149,139,142,150,150,153,153,151,143);
		wait for 10 ns;
		t_blur_matrix_int <= (144,142,147,147,141,130,122,108,144,153,153,149,139,127,118,115,151,152,154,149,144,133,121,114,155,156,148,142,134,128,124,118,154,149,149,142,136,131,122,116,150,147,147,136,132,125,120,114,150,145,141,136,132,123,109,109,146,144,140,135,128,120,114,106);
		wait for 10 ns;
		t_blur_matrix_int <= (103,109,102,96,89,91,89,85,107,111,106,99,90,97,84,85,117,112,107,99,95,93,88,91,113,110,109,102,93,94,91,86,115,116,111,105,98,96,85,94,110,115,108,103,95,88,89,94,103,112,104,100,92,85,91,92,102,103,104,97,90,86,86,92);
		wait for 10 ns;
		t_blur_matrix_int <= (101,127,168,192,214,203,178,164,97,124,161,192,213,208,183,161,99,117,154,194,211,206,188,159,95,120,151,191,210,211,191,161,96,118,143,188,214,215,195,160,97,112,146,184,208,214,199,163,100,116,135,173,206,215,203,162,96,113,129,155,200,216,204,164);
		wait for 10 ns;
		t_blur_matrix_int <= (158,143,132,122,114,106,100,98,153,152,134,120,111,106,102,100,146,139,137,129,116,105,98,94,146,140,134,130,119,107,101,96,145,136,134,130,120,113,107,96,144,139,136,125,120,114,107,96,144,144,131,129,122,114,109,100,141,135,134,123,117,122,109,102);
		wait for 10 ns;
		t_blur_matrix_int <= (93,87,85,84,77,60,34,23,95,87,87,84,79,68,35,26,90,91,91,84,81,62,32,29,89,90,90,87,82,65,26,28,94,90,90,88,77,56,27,29,96,90,92,89,74,50,27,25,93,90,89,85,76,42,31,21,95,94,90,85,68,38,23,16);
		wait for 10 ns;
		t_blur_matrix_int <= (17,19,32,26,45,30,11,63,21,25,32,32,44,22,9,57,18,30,36,34,48,22,16,44,19,31,28,40,49,23,14,41,19,29,24,37,57,23,12,32,19,28,24,35,57,16,9,28,22,21,21,33,56,15,9,21,26,19,27,40,55,15,10,16);
		wait for 10 ns;
		t_blur_matrix_int <= (141,164,134,61,37,31,16,30,137,157,138,69,34,17,12,34,137,155,141,92,33,24,17,25,134,147,132,115,26,18,12,19,128,149,111,133,29,16,12,17,128,147,113,140,38,16,20,20,130,155,118,140,62,15,9,17,119,154,119,132,85,26,11,18);
		wait for 10 ns;
		t_blur_matrix_int <= (23,18,27,25,17,23,62,102,15,24,29,21,19,27,79,112,17,24,27,17,16,41,91,116,15,26,24,15,15,52,100,114,33,24,22,21,18,70,108,120,38,26,23,16,28,79,110,115,41,31,27,20,43,96,116,114,34,29,28,20,56,105,114,113);
		wait for 10 ns;
		t_blur_matrix_int <= (118,109,110,123,139,140,138,133,113,111,109,134,140,138,136,135,113,109,118,134,141,140,136,136,115,111,121,137,142,137,138,137,116,112,131,141,144,138,135,132,113,121,135,143,140,136,134,132,112,135,153,147,140,135,136,133,110,132,153,149,136,134,134,135);
		wait for 10 ns;
		t_blur_matrix_int <= (135,132,131,128,128,131,132,130,136,131,134,131,132,133,130,131,132,134,136,130,129,130,130,131,134,136,136,131,131,133,133,129,135,136,135,132,127,130,129,128,135,133,131,133,130,127,128,129,134,138,130,133,127,130,129,128,135,131,134,129,135,127,127,128);
		wait for 10 ns;
		t_blur_matrix_int <= (130,130,130,129,128,128,130,126,135,131,130,133,129,130,129,127,128,126,137,130,128,125,125,126,130,130,129,128,128,128,126,124,129,126,127,125,129,128,128,123,129,129,126,126,128,124,128,125,125,125,125,127,128,125,124,125,125,125,127,127,125,124,123,121);
		wait for 10 ns;
		t_blur_matrix_int <= (127,125,125,122,123,120,121,120,128,124,126,125,124,121,119,117,125,125,125,123,123,121,120,116,125,129,125,120,125,124,119,116,125,124,127,123,121,121,116,114,125,121,125,124,120,120,117,113,121,124,121,120,120,115,112,110,124,124,122,122,119,115,112,108);
		wait for 10 ns;
		t_blur_matrix_int <= (116,117,115,115,112,115,139,158,119,114,114,113,115,136,156,173,115,112,112,113,129,154,171,181,115,110,112,120,148,169,179,183,111,107,114,142,162,178,184,184,110,103,128,155,175,183,188,186,105,117,144,169,180,185,186,184,110,134,161,177,183,186,186,182);
		wait for 10 ns;
		t_blur_matrix_int <= (173,181,187,188,188,187,184,182,183,187,189,189,188,185,185,182,185,188,187,187,186,185,185,182,185,185,187,185,188,186,186,184,184,183,183,186,185,184,182,184,182,182,182,184,186,184,185,185,184,185,182,186,184,186,185,186,183,181,181,184,183,185,187,192);
		wait for 10 ns;
		t_blur_matrix_int <= (182,179,178,176,178,180,180,181,181,179,178,179,182,180,181,183,182,179,179,181,183,182,184,186,184,181,182,183,185,188,191,192,184,183,186,187,190,192,193,194,186,187,190,193,196,196,196,196,192,193,195,197,198,197,198,196,196,198,200,198,198,197,195,195);
		wait for 10 ns;
		t_blur_matrix_int <= (45,47,44,44,42,46,48,39,53,44,47,46,47,46,44,43,48,49,45,47,53,47,49,40,48,48,50,45,45,43,43,38,47,50,51,43,47,39,43,44,50,49,47,47,44,46,48,45,52,48,50,45,48,47,43,38,53,57,49,49,47,45,42,39);
		wait for 10 ns;
		t_blur_matrix_int <= (39,40,31,24,24,32,62,89,39,35,29,19,18,38,66,90,33,35,30,21,20,35,57,90,38,32,25,22,14,25,59,93,38,30,22,20,16,21,58,87,32,30,21,22,11,25,56,88,29,27,24,16,10,20,54,87,37,30,25,17,11,24,59,88);
		wait for 10 ns;
		t_blur_matrix_int <= (112,126,133,147,154,153,151,150,109,124,136,140,151,150,152,150,111,121,135,146,149,152,149,149,106,125,135,146,148,151,152,150,107,124,135,146,148,152,152,156,106,123,137,143,150,152,155,152,104,123,138,145,149,154,151,153,106,122,139,146,150,152,154,153);
		wait for 10 ns;
		t_blur_matrix_int <= (153,156,157,143,133,121,108,89,158,156,158,143,135,121,107,86,153,155,154,145,136,120,110,88,151,155,155,149,136,123,108,87,154,156,154,149,138,125,108,85,154,158,156,149,141,125,110,86,154,156,159,149,141,126,108,87,157,158,157,149,140,127,108,86);
		wait for 10 ns;
		t_blur_matrix_int <= (61,45,37,46,74,105,63,63,64,39,42,38,79,103,62,57,57,40,41,38,61,119,79,83,59,42,39,38,50,81,119,106,59,42,40,42,49,62,70,80,64,44,38,44,51,59,71,92,64,43,33,45,63,91,101,83,59,44,44,70,102,100,74,70);
		wait for 10 ns;
		t_blur_matrix_int <= (71,70,83,113,134,119,76,41,81,117,141,121,107,57,16,28,134,114,82,98,102,37,23,44,89,75,83,93,89,47,32,64,89,98,98,104,99,54,24,55,83,78,96,100,89,37,41,63,71,77,81,81,59,38,45,63,72,79,83,80,55,43,38,64);
		wait for 10 ns;
		t_blur_matrix_int <= (30,60,113,84,49,103,74,25,48,100,128,69,91,66,26,25,97,109,65,83,62,34,35,31,105,78,56,75,59,84,32,51,84,63,68,61,69,34,57,66,51,56,86,72,47,58,67,46,43,73,102,55,54,55,44,35,59,98,90,50,59,43,51,31);
		wait for 10 ns;
		t_blur_matrix_int <= (26,71,43,48,31,89,122,80,36,94,61,43,52,132,112,91,64,72,101,53,84,112,87,111,73,64,104,39,97,94,91,136,51,104,78,52,90,65,101,143,50,113,36,38,88,51,102,145,93,88,20,46,108,48,94,136,116,58,19,42,112,56,71,140);
		wait for 10 ns;
		t_blur_matrix_int <= (112,39,32,33,34,25,40,22,90,68,25,29,46,31,35,18,62,113,34,35,41,27,31,19,59,114,34,19,25,33,33,19,52,74,42,15,20,20,26,21,60,48,80,13,19,29,17,28,84,31,102,21,18,21,34,47,97,23,89,39,27,43,36,21);
		wait for 10 ns;
		t_blur_matrix_int <= (24,16,20,23,13,33,53,30,14,15,14,21,17,36,58,45,11,13,12,18,27,60,90,58,11,16,14,31,30,42,81,62,17,18,18,22,52,61,54,55,28,22,18,13,33,55,38,47,24,16,8,24,38,55,79,82,19,37,9,18,30,54,106,75);
		wait for 10 ns;
		t_blur_matrix_int <= (30,27,17,32,71,113,96,41,49,21,44,51,88,142,133,55,37,18,56,73,112,162,163,87,26,50,69,93,70,157,170,109,42,118,96,83,42,56,102,73,70,120,72,51,31,79,66,28,60,108,131,99,66,60,39,15,21,38,62,84,33,18,11,10);
		wait for 10 ns;
		t_blur_matrix_int <= (80,140,125,25,15,14,14,17,32,97,130,40,7,9,5,55,20,54,107,30,6,3,12,104,15,29,55,8,5,5,43,117,17,15,25,10,15,10,82,107,14,19,22,7,27,65,100,81,9,19,8,20,104,117,102,80,12,11,6,74,149,143,138,134);
		wait for 10 ns;
		t_blur_matrix_int <= (106,96,76,109,191,190,196,201,120,86,85,152,192,196,199,131,105,88,100,175,193,198,163,22,83,88,132,192,197,190,49,14,87,98,181,197,196,92,11,15,88,131,191,153,132,23,6,12,81,122,136,140,120,36,12,11,119,125,167,156,75,10,6,19);
		wait for 10 ns;
		t_blur_matrix_int <= (66,12,12,28,36,25,38,52,15,11,10,27,43,20,29,51,10,12,10,32,48,25,32,48,13,9,11,31,57,30,36,46,13,10,10,39,66,27,38,49,13,13,9,42,74,30,36,46,12,14,18,42,74,37,37,47,17,13,12,45,78,48,33,49);
		wait for 10 ns;
		t_blur_matrix_int <= (65,74,79,87,92,90,94,97,64,74,78,85,93,91,96,95,67,69,79,86,90,92,89,93,63,73,78,92,83,90,91,97,61,71,80,84,89,92,91,95,59,68,77,82,87,89,93,95,58,73,79,82,87,89,88,95,62,74,78,88,83,93,88,92);
		wait for 10 ns;
		t_blur_matrix_int <= (106,103,113,120,120,126,125,129,98,107,109,114,119,127,126,132,100,99,108,114,119,124,123,129,99,100,106,114,111,120,118,127,98,101,107,107,113,118,118,118,99,94,99,108,113,115,120,119,95,102,103,109,108,112,120,120,95,97,103,107,109,109,112,119);
		wait for 10 ns;
		t_blur_matrix_int <= (139,142,152,148,149,149,149,142,131,135,142,148,140,145,147,144,134,128,134,142,141,144,142,143,132,127,129,132,134,140,137,140,121,127,125,125,130,137,138,133,120,119,123,130,130,131,137,131,117,121,123,124,126,131,129,131,119,120,127,126,127,127,129,133);
		wait for 10 ns;
		t_blur_matrix_int <= (145,140,137,134,124,120,106,98,145,141,136,135,128,119,103,97,141,135,134,130,123,116,106,100,135,138,139,130,121,111,103,98,133,135,128,125,114,110,99,90,135,130,127,119,114,111,96,82,133,131,125,116,108,110,82,69,129,129,125,118,114,111,86,68);
		wait for 10 ns;
		t_blur_matrix_int <= (99,98,103,95,88,89,83,88,97,98,96,94,91,82,81,87,94,95,96,90,88,84,82,85,94,92,93,91,86,82,82,84,89,86,95,99,85,84,85,78,78,89,95,99,92,87,86,84,81,96,103,100,103,103,95,86,81,98,105,100,106,107,106,89);
		wait for 10 ns;
		t_blur_matrix_int <= (99,104,128,156,195,213,209,170,92,99,129,156,193,211,214,183,88,105,125,151,180,209,219,197,89,100,121,140,169,209,220,206,90,98,121,137,161,206,223,206,93,98,115,139,157,203,223,211,89,97,108,136,161,199,224,210,81,87,108,134,163,190,212,205);
		wait for 10 ns;
		t_blur_matrix_int <= (134,134,132,126,114,115,105,102,139,141,127,124,113,112,105,98,129,131,127,122,116,112,108,97,135,136,124,123,115,113,105,100,146,129,127,122,119,113,103,103,151,118,118,120,120,111,104,97,148,116,117,117,116,107,100,94,143,116,118,116,109,104,101,92);
		wait for 10 ns;
		t_blur_matrix_int <= (96,93,91,85,63,32,23,22,96,94,89,82,52,30,14,18,94,92,90,73,47,26,20,23,95,93,83,69,44,16,16,26,94,93,83,62,30,16,20,22,91,89,85,57,18,17,21,24,93,87,77,37,20,18,20,27,89,88,66,25,15,18,19,22);
		wait for 10 ns;
		t_blur_matrix_int <= (28,28,27,42,57,13,7,12,27,37,28,40,60,11,11,17,22,35,39,44,59,15,8,15,20,35,36,45,53,13,5,16,30,38,37,43,47,21,5,14,17,33,41,45,39,26,7,13,23,35,47,42,44,24,8,12,25,35,41,44,37,23,11,18);
		wait for 10 ns;
		t_blur_matrix_int <= (107,146,117,126,94,33,12,21,95,147,115,132,103,40,10,25,78,142,129,132,112,37,6,23,68,138,139,126,118,42,10,27,56,134,139,123,120,54,18,20,45,123,141,123,129,81,23,18,27,119,145,133,132,92,24,18,19,107,147,133,124,98,35,15);
		wait for 10 ns;
		t_blur_matrix_int <= (30,29,17,21,79,111,114,113,28,23,15,42,89,117,114,111,23,20,15,53,101,117,113,112,18,22,22,68,109,117,111,116,15,18,36,83,115,115,112,117,13,14,50,95,118,119,114,121,13,16,70,105,124,120,116,127,11,16,80,114,120,121,115,134);
		wait for 10 ns;
		t_blur_matrix_int <= (120,142,140,144,138,136,138,133,122,142,140,143,141,135,137,136,131,140,141,141,136,135,132,131,130,141,140,141,137,134,123,133,138,141,137,139,135,134,130,132,143,140,138,136,133,135,134,130,142,136,136,133,133,133,131,129,140,140,136,135,136,134,129,129);
		wait for 10 ns;
		t_blur_matrix_int <= (131,136,131,129,129,126,127,127,137,134,134,132,131,130,128,130,132,134,133,130,131,131,129,130,134,135,131,132,130,131,133,129,131,131,131,134,135,132,129,127,132,130,125,127,130,130,129,128,129,133,128,129,131,129,129,134,130,129,129,130,129,128,126,127);
		wait for 10 ns;
		t_blur_matrix_int <= (127,124,125,125,124,124,123,127,124,126,126,125,124,122,122,123,127,126,128,128,126,125,123,123,125,127,129,126,123,125,124,120,129,128,131,127,124,126,124,125,129,127,128,129,126,124,124,122,130,130,127,129,126,126,132,123,131,126,128,128,125,124,124,124);
		wait for 10 ns;
		t_blur_matrix_int <= (122,119,124,119,115,115,111,111,120,119,122,117,119,115,106,111,120,118,117,120,112,111,107,124,117,117,121,115,117,110,114,137,124,115,121,116,109,110,126,157,120,118,116,112,109,115,140,169,119,117,113,108,109,122,151,178,122,113,115,106,111,136,161,181);
		wait for 10 ns;
		t_blur_matrix_int <= (123,149,172,182,185,185,183,181,138,166,180,186,187,186,183,180,152,175,183,187,185,183,181,183,167,181,185,186,184,183,182,184,176,185,187,186,184,182,182,183,183,188,186,184,186,184,184,183,185,190,187,183,183,184,185,186,187,187,186,185,183,184,184,189);
		wait for 10 ns;
		t_blur_matrix_int <= (184,181,183,184,186,189,192,196,182,182,183,187,190,194,198,199,183,184,185,191,195,198,200,202,182,185,188,195,200,202,200,202,184,190,194,199,202,203,201,200,190,194,198,203,202,202,202,197,192,195,199,202,203,200,200,197,195,198,202,200,202,200,198,196);
		wait for 10 ns;
		t_blur_matrix_int <= (199,202,202,199,197,194,195,194,203,202,202,200,197,193,194,192,202,203,203,199,196,194,194,195,203,201,201,200,200,198,196,198,201,199,200,200,201,200,198,198,197,200,200,201,201,200,201,200,198,199,199,201,202,201,201,200,199,198,202,202,201,203,200,198);
		wait for 10 ns;
		t_blur_matrix_int <= (61,51,49,54,47,50,42,40,50,53,46,48,46,44,45,42,47,48,47,44,45,45,50,40,47,53,46,45,43,46,41,39,45,51,44,48,43,40,43,41,44,51,46,43,39,48,46,42,46,51,45,46,50,49,47,42,51,48,38,42,46,46,41,40);
		wait for 10 ns;
		t_blur_matrix_int <= (34,33,31,18,12,34,62,89,34,32,32,24,18,39,69,92,35,33,35,30,30,46,78,98,37,41,38,36,34,55,83,103,32,34,40,41,47,58,88,108,35,38,41,42,52,66,92,110,40,38,35,43,58,72,94,114,38,29,28,41,63,73,96,112);
		wait for 10 ns;
		t_blur_matrix_int <= (106,122,138,145,150,149,152,150,111,122,137,145,145,151,151,152,116,125,135,143,150,152,151,154,120,128,139,145,147,151,148,154,119,129,138,142,146,146,148,149,123,132,139,145,143,147,145,150,126,131,138,144,145,147,150,151,123,132,139,140,145,147,147,152);
		wait for 10 ns;
		t_blur_matrix_int <= (152,157,159,151,143,127,106,89,153,158,156,151,141,123,110,91,153,156,157,148,144,127,108,93,154,157,157,153,142,128,108,90,151,157,160,155,144,125,112,94,154,154,159,154,144,126,111,91,151,157,156,155,143,129,111,96,155,158,160,153,144,127,114,96);
		wait for 10 ns;
		t_blur_matrix_int <= (70,62,79,80,72,62,62,64,74,59,42,44,51,56,61,68,70,47,36,46,53,58,61,64,63,46,38,50,56,60,65,69,69,44,39,48,57,57,64,65,66,50,38,47,53,58,63,63,68,49,45,48,53,58,59,65,70,47,42,47,56,62,63,67);
		wait for 10 ns;
		t_blur_matrix_int <= (68,83,88,79,53,37,38,66,67,77,85,78,52,42,44,68,68,76,80,63,49,53,48,67,73,77,87,63,61,50,53,61,73,90,83,63,50,25,46,65,75,82,81,83,26,14,36,62,67,78,104,112,36,13,37,61,73,100,121,87,44,25,38,66);
		wait for 10 ns;
		t_blur_matrix_int <= (77,91,78,55,45,18,40,84,67,108,85,54,40,10,52,139,72,112,72,50,16,16,92,109,49,65,49,39,12,65,119,80,50,52,33,9,43,108,77,42,51,39,24,31,101,71,32,30,37,45,33,102,94,39,21,30,41,64,92,108,46,31,25,30);
		wait for 10 ns;
		t_blur_matrix_int <= (101,46,26,26,97,68,51,129,72,41,46,23,87,78,62,118,38,49,64,39,73,81,66,105,36,70,70,24,75,96,70,98,60,58,50,40,69,95,53,93,58,50,52,69,82,84,67,107,49,49,49,75,97,81,89,96,44,51,42,56,80,62,88,101);
		wait for 10 ns;
		t_blur_matrix_int <= (126,29,79,98,19,28,21,21,159,52,53,126,24,23,24,45,152,78,37,132,28,20,20,52,126,117,44,134,43,9,10,20,92,145,72,120,74,7,17,28,66,126,91,120,105,19,15,25,51,102,111,120,121,57,17,30,68,81,119,89,122,89,45,42);
		wait for 10 ns;
		t_blur_matrix_int <= (27,51,10,15,27,44,31,18,33,51,11,14,17,23,36,33,36,39,29,9,13,12,16,44,19,89,100,27,19,14,6,18,14,105,139,71,13,8,9,29,16,90,140,124,19,10,11,73,22,67,102,65,30,18,43,36,51,58,70,58,39,39,37,16);
		wait for 10 ns;
		t_blur_matrix_int <= (14,27,66,82,48,14,13,14,21,103,118,19,10,15,18,19,48,118,99,22,20,21,25,19,83,98,30,12,30,27,31,32,94,63,27,13,59,57,80,79,35,37,41,51,67,79,88,128,21,47,92,84,91,101,133,165,21,59,115,110,126,146,162,171);
		wait for 10 ns;
		t_blur_matrix_int <= (17,6,8,130,147,155,155,156,11,5,28,163,160,174,166,173,9,7,82,143,150,176,173,183,37,53,94,112,132,140,153,166,89,113,78,91,91,102,172,176,161,108,77,69,89,139,207,91,141,68,75,91,118,188,149,26,72,67,57,104,172,175,46,24);
		wait for 10 ns;
		t_blur_matrix_int <= (164,167,160,90,27,10,10,17,172,157,84,22,8,6,9,16,182,104,14,11,14,13,14,19,141,40,10,7,23,22,23,15,34,15,10,14,45,62,39,17,15,16,16,18,24,36,29,23,21,28,28,24,30,34,29,27,22,33,34,30,36,37,39,35);
		wait for 10 ns;
		t_blur_matrix_int <= (17,17,9,45,77,45,34,51,22,13,11,43,74,52,40,54,20,19,8,41,87,56,43,61,19,15,19,45,90,58,41,63,15,12,22,46,95,69,46,58,22,15,13,50,97,65,45,57,24,19,19,50,95,72,47,61,24,20,25,47,89,77,56,64);
		wait for 10 ns;
		t_blur_matrix_int <= (59,75,79,87,87,91,86,91,60,75,79,82,82,87,91,89,66,70,76,84,82,86,90,92,67,77,74,84,85,84,90,90,71,74,79,82,85,86,88,94,71,75,80,83,84,85,89,90,71,76,83,83,85,89,83,89,72,79,86,86,87,90,92,93);
		wait for 10 ns;
		t_blur_matrix_int <= (94,97,107,102,109,107,114,118,94,101,100,102,108,106,121,112,92,99,99,106,112,110,110,119,93,98,98,105,108,112,111,116,90,95,97,99,109,110,109,115,87,94,96,96,103,106,111,110,93,96,98,102,104,108,108,108,93,96,103,103,103,104,102,108);
		wait for 10 ns;
		t_blur_matrix_int <= (117,117,115,121,126,122,129,127,119,119,123,120,122,126,127,128,117,114,118,117,127,126,128,127,117,111,119,119,122,122,122,127,111,112,118,117,125,117,122,127,111,114,115,114,122,123,123,122,111,106,112,117,120,121,126,127,105,110,114,121,121,121,121,123);
		wait for 10 ns;
		t_blur_matrix_int <= (129,128,126,118,112,110,83,70,130,127,130,120,114,106,97,79,128,128,129,120,117,116,102,80,131,126,131,125,116,118,111,93,128,128,128,127,120,119,115,108,129,128,130,126,125,124,121,115,130,129,128,128,124,128,120,117,125,128,127,126,121,121,122,120);
		wait for 10 ns;
		t_blur_matrix_int <= (86,99,97,94,85,97,96,91,94,97,86,30,18,36,61,66,86,91,80,55,46,66,66,55,81,85,89,91,90,93,91,78,102,95,84,87,90,93,96,81,109,107,96,96,96,106,123,116,117,112,108,105,108,125,155,158,116,116,112,112,123,140,177,180);
		wait for 10 ns;
		t_blur_matrix_int <= (79,80,96,118,152,183,194,189,81,83,86,97,138,173,186,152,53,72,81,91,118,161,173,144,75,70,81,90,122,169,158,144,81,101,134,157,171,171,153,139,111,138,177,185,180,172,151,140,123,145,179,181,179,174,154,134,143,152,180,183,180,176,150,132);
		wait for 10 ns;
		t_blur_matrix_int <= (127,117,116,114,112,109,104,95,123,119,116,116,111,104,94,92,137,116,116,112,106,105,100,96,131,123,116,109,105,101,95,95,128,122,117,108,103,98,98,88,123,121,115,112,102,101,94,76,125,117,112,107,98,97,94,57,118,113,115,105,103,102,84,27);
		wait for 10 ns;
		t_blur_matrix_int <= (91,81,38,17,17,20,22,27,90,65,22,17,20,21,27,31,86,38,22,20,21,21,26,23,70,25,21,30,26,19,29,27,46,19,22,26,24,24,29,27,28,23,20,26,23,22,31,32,26,28,22,23,20,26,29,37,24,27,25,26,25,27,41,38);
		wait for 10 ns;
		t_blur_matrix_int <= (24,30,47,33,39,16,16,15,30,37,48,29,40,19,22,12,28,38,41,38,41,19,23,19,32,43,44,38,44,16,22,22,30,56,48,41,41,19,22,16,37,62,46,52,36,26,37,17,32,70,37,57,37,24,39,19,37,64,38,49,34,31,36,29);
		wait for 10 ns;
		t_blur_matrix_int <= (13,94,146,146,120,100,35,19,10,87,139,146,109,111,49,20,8,63,141,149,102,121,51,14,7,44,136,145,112,126,64,14,10,30,131,152,107,124,71,23,12,21,118,153,106,116,68,26,13,13,105,152,106,118,60,39,15,16,86,152,119,119,62,54);
		wait for 10 ns;
		t_blur_matrix_int <= (12,22,86,122,125,117,122,139,19,45,99,126,123,119,126,140,31,60,109,125,120,118,129,137,34,79,119,125,122,123,132,140,35,96,121,122,119,123,138,139,45,108,123,121,123,128,140,137,65,113,122,119,119,131,140,134,85,118,124,117,124,130,140,134);
		wait for 10 ns;
		t_blur_matrix_int <= (141,139,136,133,131,133,132,128,138,137,134,135,135,132,128,130,138,135,133,133,131,130,130,129,139,138,135,134,131,129,129,129,138,134,133,134,131,131,132,129,134,136,136,133,129,131,132,130,134,133,136,135,130,132,132,128,137,136,134,131,130,130,130,131);
		wait for 10 ns;
		t_blur_matrix_int <= (133,131,130,130,134,131,132,128,130,127,128,129,127,129,124,123,128,129,127,133,129,128,127,126,130,129,133,130,126,129,127,129,127,127,130,130,130,128,128,127,130,128,126,129,130,130,127,126,128,128,126,127,128,129,127,124,128,128,128,129,128,123,125,126);
		wait for 10 ns;
		t_blur_matrix_int <= (127,131,127,129,126,127,124,119,125,130,125,123,123,122,125,121,126,124,124,123,124,127,122,119,127,125,127,124,125,121,121,121,124,127,126,124,121,122,121,123,127,126,125,125,127,120,120,118,125,125,128,125,123,124,121,121,127,126,127,125,126,118,119,120);
		wait for 10 ns;
		t_blur_matrix_int <= (118,116,112,108,116,149,169,183,120,112,112,107,124,153,173,183,119,115,111,112,131,161,180,185,118,114,109,116,141,165,183,186,116,112,110,121,148,173,184,187,115,114,111,124,155,177,186,183,112,113,111,133,156,176,185,186,114,109,114,136,165,181,187,185);
		wait for 10 ns;
		t_blur_matrix_int <= (187,185,183,182,182,185,189,194,187,187,186,185,186,189,194,197,188,187,186,186,188,191,197,198,186,186,187,186,190,195,201,199,187,184,186,190,195,196,201,202,187,186,188,191,196,199,202,200,185,186,189,194,198,201,202,200,186,188,193,198,201,203,202,200);
		wait for 10 ns;
		t_blur_matrix_int <= (196,198,198,200,199,198,201,200,198,199,197,198,199,200,203,202,199,199,198,199,200,200,203,205,201,201,201,202,201,200,203,205,199,200,200,200,200,202,205,205,200,199,199,199,199,202,204,203,200,198,198,200,201,202,203,204,200,198,198,200,201,202,202,203);
		wait for 10 ns;
		t_blur_matrix_int <= (199,200,201,204,203,202,201,199,203,203,203,203,205,203,201,199,203,203,204,204,205,202,200,201,204,203,203,204,202,201,199,200,204,203,205,203,200,200,200,202,204,204,206,202,202,200,203,204,204,205,203,203,203,205,205,204,203,205,203,208,203,206,204,204);
		wait for 10 ns;
		t_blur_matrix_int <= (41,46,36,42,40,39,41,42,43,44,37,42,40,39,42,35,44,40,40,39,38,31,37,38,41,36,37,36,35,38,36,37,43,32,31,32,34,41,38,36,40,28,29,30,34,35,38,36,28,28,28,28,28,31,37,36,29,27,27,30,33,35,37,31);
		wait for 10 ns;
		t_blur_matrix_int <= (33,30,29,40,55,79,99,114,31,30,30,40,62,77,98,112,34,33,36,44,53,73,93,112,28,33,38,44,53,71,91,109,32,31,34,38,52,68,93,109,35,28,33,44,50,69,96,111,33,28,31,42,51,67,95,112,29,27,38,46,57,75,98,118);
		wait for 10 ns;
		t_blur_matrix_int <= (125,134,137,145,145,147,146,149,124,133,140,140,148,145,144,152,123,129,139,141,146,149,149,153,123,132,138,144,147,147,152,153,126,131,140,146,148,150,150,154,125,138,138,144,149,149,149,152,127,139,144,147,151,150,155,155,125,135,141,152,154,156,155,158);
		wait for 10 ns;
		t_blur_matrix_int <= (153,159,156,151,145,129,113,92,153,159,159,155,145,132,113,96,151,156,158,155,143,134,116,92,155,157,160,158,148,131,117,94,156,160,161,155,149,130,114,94,154,161,160,156,148,134,116,89,158,160,157,158,146,130,115,90,157,160,158,155,147,131,110,89);
		wait for 10 ns;
		t_blur_matrix_int <= (68,51,42,47,50,53,60,59,71,49,36,42,52,52,59,80,67,46,38,46,52,48,65,108,71,44,34,45,49,59,103,104,73,41,37,39,47,90,109,67,67,45,38,41,65,114,73,58,68,41,33,54,105,88,54,56,67,45,38,110,102,58,48,58);
		wait for 10 ns;
		t_blur_matrix_int <= (89,118,90,80,47,38,41,49,120,86,85,81,30,34,43,60,90,75,97,78,31,33,63,84,71,70,100,71,32,53,61,77,64,72,92,62,37,42,23,88,61,73,108,61,32,16,35,89,71,97,114,51,24,18,52,32,101,121,108,49,26,40,60,17);
		wait for 10 ns;
		t_blur_matrix_int <= (71,110,79,41,39,21,28,24,107,89,17,22,65,29,32,28,108,60,18,27,45,52,43,40,92,39,25,28,35,50,41,50,72,31,34,29,51,39,36,58,97,33,36,32,43,36,32,43,70,41,38,36,45,41,33,29,29,31,42,39,49,44,37,28);
		wait for 10 ns;
		t_blur_matrix_int <= (48,47,47,45,59,46,87,82,45,40,48,40,57,46,65,97,45,29,65,44,47,45,47,93,42,46,55,54,41,45,44,75,43,69,56,64,52,46,54,54,40,58,83,65,74,62,60,51,33,65,107,69,81,77,62,51,30,73,122,97,84,74,86,65);
		wait for 10 ns;
		t_blur_matrix_int <= (73,54,108,80,132,99,50,50,42,57,96,101,128,103,65,36,34,51,92,109,96,99,98,70,67,26,36,92,120,90,116,120,70,64,27,43,107,98,115,132,42,90,59,29,47,67,99,115,43,47,91,60,53,79,75,102,61,38,53,93,102,78,41,77);
		wait for 10 ns;
		t_blur_matrix_int <= (74,63,60,55,22,27,31,16,110,61,32,29,17,11,32,52,137,25,26,12,36,43,59,78,91,7,19,13,48,98,95,75,48,16,16,47,97,114,150,149,104,32,20,84,66,94,151,191,78,85,93,136,107,104,162,182,51,47,105,111,93,139,178,187);
		wait for 10 ns;
		t_blur_matrix_int <= (42,142,136,132,149,161,174,128,79,122,127,135,161,182,173,73,73,100,131,144,172,185,99,67,80,111,141,155,187,131,68,57,126,148,179,184,157,61,74,66,189,193,188,163,69,75,55,80,200,197,179,83,75,66,67,123,203,192,120,60,74,65,99,181);
		wait for 10 ns;
		t_blur_matrix_int <= (61,62,64,107,185,57,16,17,71,59,81,162,94,17,14,18,59,65,136,129,23,15,23,22,63,108,160,23,16,13,34,42,94,162,64,22,18,16,50,59,146,113,13,16,14,16,43,64,165,24,18,15,21,16,24,51,73,13,20,24,25,15,21,45);
		wait for 10 ns;
		t_blur_matrix_int <= (20,21,23,20,22,29,40,36,29,21,20,16,21,23,45,30,29,27,21,23,18,31,43,39,25,24,17,24,24,25,44,44,26,23,15,26,22,26,39,55,18,21,14,26,25,29,45,44,17,17,17,22,25,38,37,40,29,12,18,19,27,31,30,43);
		wait for 10 ns;
		t_blur_matrix_int <= (24,17,17,30,89,78,57,63,21,23,8,31,81,75,70,60,22,20,16,22,74,71,80,49,27,18,10,19,80,66,76,47,34,15,13,18,70,62,76,52,33,19,11,22,73,55,72,46,43,14,14,17,81,51,67,44,50,12,11,17,71,39,68,51);
		wait for 10 ns;
		t_blur_matrix_int <= (73,75,83,83,87,87,88,87,70,74,80,81,86,88,94,92,71,73,79,82,86,91,88,91,60,72,74,86,84,87,89,90,56,69,74,79,86,88,89,93,51,63,74,84,83,89,92,93,49,59,71,77,83,91,95,88,41,59,69,82,79,93,94,89);
		wait for 10 ns;
		t_blur_matrix_int <= (94,94,100,101,106,107,103,102,87,97,99,98,104,100,104,103,90,93,101,97,103,108,100,100,92,94,100,100,104,108,102,106,91,92,101,100,100,103,104,103,88,93,95,95,98,101,106,106,88,88,91,95,95,99,103,108,91,87,93,94,99,103,102,105);
		wait for 10 ns;
		t_blur_matrix_int <= (104,103,108,113,117,118,120,120,108,105,107,108,112,115,116,118,107,99,106,103,104,111,114,115,100,99,102,102,107,105,107,111,102,99,100,104,109,106,101,106,101,103,101,106,99,96,92,91,107,106,106,114,91,57,53,70,108,110,111,110,84,58,59,46);
		wait for 10 ns;
		t_blur_matrix_int <= (117,122,121,126,121,118,119,119,115,121,121,127,122,115,114,121,112,113,115,124,114,119,113,117,112,112,110,115,110,112,113,114,110,103,102,112,113,112,105,110,95,100,101,110,105,111,108,110,83,88,94,95,92,91,87,82,41,47,53,57,58,64,72,62);
		wait for 10 ns;
		t_blur_matrix_int <= (116,116,118,121,127,154,190,186,122,120,122,123,136,164,197,192,120,125,127,129,141,166,199,193,117,122,123,130,140,169,193,199,120,128,134,129,132,132,147,154,106,104,100,97,93,90,106,104,78,79,80,74,75,73,81,87,59,56,52,47,52,62,71,76);
		wait for 10 ns;
		t_blur_matrix_int <= (158,152,184,187,185,179,146,130,167,152,187,191,181,174,150,131,166,149,174,193,184,174,146,122,175,168,195,191,184,176,150,115,179,181,155,138,136,153,145,102,118,122,111,102,104,116,105,76,101,97,62,51,67,78,61,70,81,68,62,54,68,86,81,92);
		wait for 10 ns;
		t_blur_matrix_int <= (120,111,114,103,101,96,55,20,113,114,111,104,104,88,27,22,109,112,107,106,100,64,22,22,106,105,106,105,97,30,18,20,94,100,108,105,68,25,20,18,91,107,111,100,31,24,19,23,97,112,111,75,23,22,20,23,107,116,104,36,19,22,18,24);
		wait for 10 ns;
		t_blur_matrix_int <= (26,27,21,22,22,24,40,35,21,24,24,25,20,30,40,37,23,25,23,23,27,28,38,36,21,37,27,23,24,33,36,41,26,38,25,21,29,27,42,41,28,24,26,27,30,29,43,39,29,23,22,22,29,30,51,27,28,20,22,28,26,42,42,31);
		wait for 10 ns;
		t_blur_matrix_int <= (43,58,36,49,32,32,28,17,48,54,38,46,30,38,25,21,51,53,42,48,23,36,29,22,49,48,37,46,32,34,32,18,51,56,39,48,44,34,40,17,49,53,43,52,38,30,38,19,49,44,41,56,37,21,37,28,56,42,48,54,34,13,47,41);
		wait for 10 ns;
		t_blur_matrix_int <= (11,10,64,145,129,117,58,78,12,11,61,135,123,109,61,86,13,13,63,127,137,104,62,99,13,9,55,120,138,106,69,96,10,8,41,118,145,100,80,105,10,12,28,117,143,89,90,106,11,11,23,103,141,88,106,111,16,17,21,90,139,105,118,109);
		wait for 10 ns;
		t_blur_matrix_int <= (93,119,122,114,126,136,137,133,98,118,122,117,127,136,134,133,106,116,119,123,128,137,131,137,108,114,118,125,135,138,134,133,113,116,119,122,132,136,135,135,116,122,118,122,135,137,135,136,121,119,124,118,134,137,136,137,124,120,123,125,138,134,145,133);
		wait for 10 ns;
		t_blur_matrix_int <= (134,133,132,131,129,130,130,127,135,135,131,131,129,128,126,128,135,130,135,133,133,127,129,131,136,136,129,132,129,127,125,127,134,133,130,130,131,128,125,128,134,131,129,129,129,125,127,123,130,131,134,130,129,130,128,126,133,133,134,132,130,131,127,128);
		wait for 10 ns;
		t_blur_matrix_int <= (129,127,127,126,123,125,124,126,126,129,131,129,128,122,124,126,127,126,128,128,125,126,125,126,127,126,131,126,126,128,125,123,130,134,127,129,126,127,120,125,127,132,127,127,130,129,125,124,131,128,129,127,130,126,126,125,126,130,129,125,126,129,126,125);
		wait for 10 ns;
		t_blur_matrix_int <= (125,125,124,129,124,119,122,120,120,125,125,125,125,122,119,119,125,127,125,125,120,122,115,112,125,124,123,122,123,119,116,114,125,124,123,122,122,117,117,115,126,124,121,123,118,120,116,114,126,124,123,122,124,121,116,114,123,123,125,123,122,120,116,110);
		wait for 10 ns;
		t_blur_matrix_int <= (114,110,116,144,166,183,185,188,114,108,116,145,172,184,186,184,109,109,119,151,174,184,187,186,111,107,122,152,174,186,186,189,109,106,122,156,174,186,189,195,108,104,126,155,176,185,193,196,107,103,131,158,176,190,196,201,106,106,132,165,179,189,199,202);
		wait for 10 ns;
		t_blur_matrix_int <= (186,191,197,200,203,202,201,198,188,195,199,203,202,201,200,199,191,197,200,203,202,201,201,200,196,200,203,202,202,200,201,201,196,202,206,203,203,200,201,202,200,205,204,203,201,201,202,202,203,205,203,204,204,203,203,201,206,204,205,203,205,202,202,200);
		wait for 10 ns;
		t_blur_matrix_int <= (200,199,199,200,203,202,201,203,200,202,200,201,203,200,201,204,200,202,201,201,202,200,202,203,203,202,202,199,200,202,206,207,203,203,204,202,202,203,205,204,202,204,202,202,204,204,207,206,201,202,201,202,205,205,208,207,202,202,204,204,204,204,206,206);
		wait for 10 ns;
		t_blur_matrix_int <= (204,206,205,205,205,206,204,205,204,205,205,204,205,204,203,206,208,206,205,203,205,206,206,206,207,205,207,206,204,205,205,206,210,208,207,206,205,207,206,205,207,209,208,207,206,208,206,206,207,208,208,206,206,207,207,210,207,210,211,208,207,208,208,206);
		wait for 10 ns;
		t_blur_matrix_int <= (25,28,27,28,29,31,37,32,29,28,30,28,30,29,31,31,27,30,28,30,31,32,36,34,29,29,24,27,30,30,29,31,31,24,26,28,26,22,28,27,21,21,24,25,25,24,25,25,37,25,20,22,22,32,27,25,26,22,25,28,20,22,21,17);
		wait for 10 ns;
		t_blur_matrix_int <= (30,32,35,56,58,75,96,117,28,34,43,61,66,80,100,115,25,30,43,55,63,75,96,115,25,27,47,58,64,71,94,113,24,26,43,56,63,66,93,111,23,28,47,56,68,64,89,110,27,27,51,65,54,61,86,105,22,33,60,66,61,60,86,104);
		wait for 10 ns;
		t_blur_matrix_int <= (125,137,144,151,152,155,156,155,125,136,143,152,156,154,156,158,125,133,139,151,153,156,158,159,125,134,140,147,154,157,159,158,125,133,140,150,152,159,159,160,121,131,137,146,157,159,157,162,119,128,134,149,157,161,158,159,114,124,131,147,155,157,159,158);
		wait for 10 ns;
		t_blur_matrix_int <= (156,161,162,155,143,130,110,90,162,162,161,153,143,129,113,86,161,163,161,156,144,132,111,86,161,161,158,153,142,144,125,107,162,163,163,154,146,141,148,110,161,160,163,155,145,130,116,89,156,163,161,155,145,128,113,91,161,162,165,152,143,131,113,91);
		wait for 10 ns;
		t_blur_matrix_int <= (66,47,91,113,66,45,50,75,67,103,124,65,42,46,59,97,104,123,70,41,45,47,75,117,111,67,36,36,43,57,96,120,77,38,31,36,48,81,129,81,64,40,34,40,59,122,103,68,64,41,33,37,84,127,69,66,65,40,29,39,89,117,63,70);
		wait for 10 ns;
		t_blur_matrix_int <= (113,109,94,43,27,50,35,25,113,90,80,56,39,38,45,25,86,79,74,57,41,34,84,39,73,72,69,43,49,50,120,41,67,79,60,28,38,84,102,32,72,87,56,29,26,116,93,18,76,78,35,28,38,125,83,14,81,55,24,30,50,116,62,21);
		wait for 10 ns;
		t_blur_matrix_int <= (16,37,43,44,52,36,48,41,29,20,28,24,56,36,40,56,32,14,20,20,66,43,32,74,15,17,15,37,77,42,33,70,23,24,20,46,76,32,64,57,21,26,24,69,68,26,58,55,23,18,23,80,48,24,33,60,22,20,39,72,38,29,21,38);
		wait for 10 ns;
		t_blur_matrix_int <= (32,71,118,108,76,72,74,78,25,82,149,103,48,70,75,75,23,87,156,101,42,40,72,87,34,101,154,101,49,31,61,60,53,130,130,94,97,31,57,70,58,154,104,68,121,68,67,100,69,175,117,48,81,113,86,108,102,167,127,71,52,130,97,110);
		wait for 10 ns;
		t_blur_matrix_int <= (85,68,59,76,124,73,38,50,79,80,70,72,50,67,67,57,94,67,60,65,38,45,86,80,75,101,80,63,52,45,64,73,37,78,105,83,83,75,90,80,52,41,70,109,78,119,111,84,61,43,35,79,127,113,78,111,71,59,54,91,109,119,99,77);
		wait for 10 ns;
		t_blur_matrix_int <= (33,62,103,109,98,97,187,215,75,94,125,109,95,87,143,216,102,104,122,111,98,79,120,203,119,113,123,107,86,104,175,176,129,131,119,115,72,127,203,112,101,143,128,112,75,126,187,104,62,118,94,122,84,144,194,130,55,102,77,99,81,169,172,123);
		wait for 10 ns;
		t_blur_matrix_int <= (205,172,75,69,56,92,168,125,188,112,71,69,87,146,166,35,132,69,79,103,154,173,69,27,63,87,106,152,149,94,21,29,82,116,144,185,105,30,31,28,119,144,183,122,44,28,32,30,151,165,165,41,30,28,28,32,155,174,55,23,26,30,29,26);
		wait for 10 ns;
		t_blur_matrix_int <= (22,20,23,21,21,20,17,35,23,27,28,26,23,17,22,34,30,28,28,26,21,18,17,25,20,27,27,29,24,19,16,18,26,29,34,33,29,22,21,29,28,30,34,28,42,29,28,30,32,30,30,32,28,21,26,32,25,28,32,31,30,20,21,29);
		wait for 10 ns;
		t_blur_matrix_int <= (32,20,18,25,26,31,27,39,31,16,21,27,33,32,29,34,27,23,15,21,33,26,33,33,27,28,22,19,26,31,32,34,27,24,28,22,26,40,28,35,28,21,33,31,33,30,39,35,25,24,28,33,35,30,38,33,22,24,33,28,32,31,30,31);
		wait for 10 ns;
		t_blur_matrix_int <= (52,21,17,17,70,42,61,54,49,28,18,22,66,41,54,53,43,31,17,25,58,35,56,55,44,39,18,23,42,33,55,54,42,40,19,27,54,46,55,49,44,43,31,21,45,48,50,50,39,39,28,24,36,49,45,54,30,35,27,25,29,45,36,58);
		wait for 10 ns;
		t_blur_matrix_int <= (46,54,64,76,83,84,91,86,49,53,63,77,79,83,89,83,37,47,57,73,74,75,84,79,34,51,59,66,73,76,82,80,33,42,54,66,71,75,76,77,34,43,45,59,66,68,67,75,31,39,39,49,62,70,69,66,35,35,43,45,52,60,64,67);
		wait for 10 ns;
		t_blur_matrix_int <= (84,89,92,93,98,98,97,100,83,88,89,88,94,97,100,102,83,86,86,90,89,91,94,103,80,85,84,83,88,93,90,97,76,82,82,89,88,95,89,95,79,82,85,88,88,96,98,97,74,77,80,82,84,90,91,92,71,68,78,79,84,87,92,92);
		wait for 10 ns;
		t_blur_matrix_int <= (115,112,112,110,91,86,88,82,112,115,113,109,109,103,90,86,109,111,110,110,115,103,96,92,108,106,108,115,112,109,103,98,103,104,105,109,112,109,104,99,99,101,102,104,104,107,108,99,99,96,102,100,107,106,102,104,95,96,104,102,105,108,103,102);
		wait for 10 ns;
		t_blur_matrix_int <= (69,61,59,63,69,75,79,77,86,84,81,78,75,84,89,96,86,87,84,86,75,76,81,89,88,87,82,85,86,89,81,81,96,93,87,84,85,88,89,84,98,94,95,89,91,87,80,81,99,96,95,91,94,90,88,84,98,99,96,93,96,92,97,99);
		wait for 10 ns;
		t_blur_matrix_int <= (79,78,75,77,78,75,85,95,89,109,117,123,132,132,145,160,101,120,140,154,155,154,158,168,91,106,109,117,124,120,110,111,83,94,99,96,107,104,99,98,81,88,89,94,100,92,91,86,81,78,77,81,79,77,79,84,95,90,87,90,94,97,104,117);
		wait for 10 ns;
		t_blur_matrix_int <= (101,106,99,86,92,107,102,105,165,158,118,95,98,112,117,109,175,160,110,96,104,118,119,108,122,119,95,107,113,120,116,109,98,95,102,115,117,122,108,100,86,99,117,121,114,115,105,67,102,126,121,110,113,113,75,41,122,124,111,104,111,106,32,41);
		wait for 10 ns;
		t_blur_matrix_int <= (113,110,67,20,22,23,22,29,112,95,29,19,23,22,22,26,105,53,19,18,19,23,24,26,87,20,19,19,18,21,30,20,52,20,24,24,21,26,28,22,35,12,24,21,26,28,22,27,27,19,19,15,18,24,18,28,24,20,23,21,18,28,28,27);
		wait for 10 ns;
		t_blur_matrix_int <= (25,22,22,27,27,45,30,31,22,23,21,29,32,37,27,38,18,14,23,28,26,22,23,44,19,16,21,24,39,19,19,43,25,18,28,22,34,22,22,46,30,25,26,28,33,21,22,52,31,33,23,25,29,20,23,67,42,36,31,27,27,25,22,71);
		wait for 10 ns;
		t_blur_matrix_int <= (53,46,42,55,33,19,46,50,57,45,45,53,40,24,43,54,63,40,49,47,24,25,40,60,66,44,57,52,35,36,35,63,56,37,55,49,39,39,28,67,56,39,56,47,47,32,28,71,50,47,53,51,45,31,35,59,50,45,55,59,39,30,36,61);
		wait for 10 ns;
		t_blur_matrix_int <= (17,17,19,76,136,109,126,113,19,18,19,66,139,119,125,114,19,16,18,62,144,127,124,120,23,21,24,61,139,131,122,126,21,21,22,62,134,136,126,126,24,26,21,59,133,142,124,128,25,23,25,56,126,145,123,128,30,34,24,51,132,150,126,133);
		wait for 10 ns;
		t_blur_matrix_int <= (125,120,126,125,136,137,136,135,129,119,127,128,140,137,136,132,128,120,127,129,138,138,137,139,134,121,129,129,137,139,139,138,134,123,130,133,137,138,137,136,133,127,130,137,139,138,135,137,130,123,131,136,138,135,135,136,127,124,133,136,138,139,135,139);
		wait for 10 ns;
		t_blur_matrix_int <= (131,133,132,133,131,130,134,128,131,134,135,131,135,130,132,128,132,135,132,132,131,135,133,131,138,140,135,134,134,132,133,135,132,134,137,133,133,132,136,132,136,134,136,138,136,134,133,132,132,136,135,134,136,134,133,138,135,137,135,136,135,136,138,138);
		wait for 10 ns;
		t_blur_matrix_int <= (127,129,126,129,132,130,126,126,128,128,125,125,127,127,127,122,132,130,130,126,132,126,125,125,130,132,131,133,128,123,125,125,133,129,129,135,128,127,125,129,131,133,131,129,130,127,126,126,135,132,131,132,130,131,126,127,138,134,133,134,130,129,127,127);
		wait for 10 ns;
		t_blur_matrix_int <= (124,125,125,124,124,118,117,111,127,126,123,125,122,118,117,109,129,127,123,125,122,123,111,111,128,125,121,126,120,118,115,107,127,126,126,122,126,119,114,110,126,124,121,118,120,116,112,108,125,124,121,123,120,117,111,104,126,125,123,122,121,113,111,104);
		wait for 10 ns;
		t_blur_matrix_int <= (106,109,139,167,184,195,201,204,102,109,137,170,187,196,206,205,102,110,143,173,192,203,206,208,103,109,144,178,195,205,209,208,100,110,145,184,202,206,210,210,100,107,148,186,201,209,211,210,95,106,150,188,205,212,212,209,95,103,148,189,206,212,213,210);
		wait for 10 ns;
		t_blur_matrix_int <= (206,205,204,205,204,203,204,201,207,206,204,204,206,205,206,203,205,205,206,203,205,205,205,204,206,205,206,203,206,206,207,206,208,206,207,204,206,206,208,208,208,206,207,207,207,207,209,210,208,207,207,207,208,210,211,211,208,209,209,209,208,210,211,211);
		wait for 10 ns;
		t_blur_matrix_int <= (203,204,205,204,205,205,206,207,206,206,206,206,208,209,209,208,205,205,206,206,207,207,209,209,208,206,207,208,209,208,208,207,209,208,209,210,211,209,206,203,210,210,210,209,207,204,202,199,213,211,208,205,204,201,200,198,209,207,205,203,202,200,200,201);
		wait for 10 ns;
		t_blur_matrix_int <= (208,209,209,208,207,207,207,205,208,207,206,206,206,206,206,205,208,207,206,206,204,205,205,202,206,203,202,204,201,200,201,200,204,202,199,200,200,198,197,198,198,198,197,197,198,199,198,197,199,198,199,201,200,201,203,202,202,203,204,204,203,204,205,204);
		wait for 10 ns;
		t_blur_matrix_int <= (28,21,24,23,22,21,22,21,28,25,24,24,21,18,18,19,21,22,21,22,22,23,22,23,17,22,20,23,23,21,24,26,20,23,20,22,21,18,24,21,21,20,28,26,17,17,25,23,24,17,26,28,23,21,22,20,24,23,19,20,20,14,22,27);
		wait for 10 ns;
		t_blur_matrix_int <= (17,44,75,70,69,73,87,100,19,51,73,75,70,73,91,103,29,60,70,72,69,74,92,100,28,54,75,75,68,75,93,100,31,59,72,74,70,70,92,103,35,53,60,65,65,72,92,103,27,45,56,66,71,80,96,104,25,35,53,67,71,83,99,99);
		wait for 10 ns;
		t_blur_matrix_int <= (112,122,132,146,154,156,157,158,111,118,130,144,151,157,155,157,113,118,131,147,150,154,157,155,110,124,132,142,155,153,154,157,109,120,135,143,154,158,155,158,108,124,133,146,153,155,155,153,110,124,134,146,152,155,153,156,113,123,134,146,151,151,151,155);
		wait for 10 ns;
		t_blur_matrix_int <= (156,159,162,154,146,131,117,94,157,158,160,153,145,136,116,95,155,158,158,151,140,129,115,93,157,157,157,156,142,133,113,91,157,155,159,153,143,132,115,92,157,158,159,154,144,134,114,93,157,157,160,154,146,133,112,95,154,159,157,154,146,134,117,93);
		wait for 10 ns;
		t_blur_matrix_int <= (66,41,29,35,88,112,60,66,67,43,31,37,69,105,71,72,67,49,35,37,58,92,82,77,65,46,30,43,56,76,72,73,66,43,30,44,52,78,72,75,69,42,33,44,56,70,79,47,64,42,32,40,52,69,80,29,65,41,31,37,51,91,50,32);
		wait for 10 ns;
		t_blur_matrix_int <= (57,49,39,31,51,97,32,27,67,53,38,55,51,67,30,26,51,45,44,74,62,56,29,21,56,46,52,59,70,50,33,27,38,40,43,34,92,47,29,30,34,36,32,38,107,41,33,35,26,30,25,46,93,60,25,36,21,25,40,61,61,52,24,38);
		wait for 10 ns;
		t_blur_matrix_int <= (22,14,45,63,29,40,25,27,21,17,51,60,26,41,31,33,15,19,57,58,19,31,34,26,18,18,62,54,22,25,34,41,25,19,61,50,19,33,31,50,28,25,51,50,22,32,24,44,41,23,49,42,20,29,18,23,40,34,46,44,23,26,26,17);
		wait for 10 ns;
		t_blur_matrix_int <= (128,150,123,112,59,102,123,111,106,148,112,78,109,77,146,112,87,120,89,85,95,83,113,124,79,113,80,65,88,100,93,115,76,100,88,36,38,51,96,104,93,105,87,38,32,30,54,89,92,115,115,50,28,43,55,73,82,130,115,79,29,56,53,67);
		wait for 10 ns;
		t_blur_matrix_int <= (84,83,107,74,65,107,105,67,87,97,89,49,69,98,109,68,92,94,78,59,57,66,110,79,103,108,95,83,57,52,121,82,122,114,106,102,79,56,123,97,118,115,89,114,114,87,103,109,87,101,106,122,120,90,95,99,87,75,101,97,134,130,125,94);
		wait for 10 ns;
		t_blur_matrix_int <= (45,109,100,95,86,159,184,166,38,96,81,102,101,189,202,190,69,108,58,90,72,149,199,138,76,112,54,75,80,117,185,58,71,129,65,52,85,88,172,40,101,119,71,69,73,64,47,42,116,125,76,69,71,79,37,43,114,130,141,51,66,76,73,34);
		wait for 10 ns;
		t_blur_matrix_int <= (191,81,30,28,26,27,25,26,116,36,20,21,27,32,22,24,35,27,25,27,29,33,31,28,31,32,24,23,27,23,26,26,57,31,25,28,30,30,24,30,55,30,30,27,36,24,24,30,35,34,24,27,28,28,22,25,32,32,29,30,28,30,30,29);
		wait for 10 ns;
		t_blur_matrix_int <= (23,33,29,31,33,23,26,33,23,28,28,32,29,19,22,33,26,26,32,31,27,21,25,34,18,34,39,28,26,18,24,33,22,44,36,30,27,15,28,33,25,34,33,34,25,21,27,38,23,31,31,35,23,22,29,40,32,37,42,44,27,20,28,40);
		wait for 10 ns;
		t_blur_matrix_int <= (26,29,28,26,34,30,30,31,20,27,28,22,25,30,34,30,25,26,30,20,18,20,32,30,21,24,28,20,20,22,23,29,23,18,29,28,20,21,23,23,23,27,24,31,19,20,22,24,22,24,24,35,29,18,24,20,23,27,31,27,31,23,25,28);
		wait for 10 ns;
		t_blur_matrix_int <= (32,34,39,25,24,36,31,51,31,36,35,23,21,32,32,36,28,33,37,23,20,29,35,32,25,28,33,29,24,25,34,31,28,30,27,29,28,27,33,29,32,30,28,25,28,28,36,28,23,32,32,26,33,24,28,34,24,25,33,31,37,38,26,30);
		wait for 10 ns;
		t_blur_matrix_int <= (38,29,43,43,53,54,60,68,43,28,35,38,37,52,53,65,44,25,29,42,30,34,48,60,34,25,28,47,34,18,30,45,37,34,24,44,43,19,18,25,34,39,26,41,43,26,17,15,33,40,26,34,42,42,23,19,32,35,29,34,45,42,33,23);
		wait for 10 ns;
		t_blur_matrix_int <= (68,73,74,82,86,90,89,92,67,70,72,75,83,90,85,93,61,66,70,73,77,87,91,92,49,59,64,65,74,81,85,95,38,48,60,59,66,75,86,89,19,35,44,47,56,70,79,85,17,17,29,40,48,62,73,82,21,18,21,25,44,45,56,60);
		wait for 10 ns;
		t_blur_matrix_int <= (97,95,98,105,101,102,101,101,97,99,105,99,101,102,106,105,95,100,104,100,104,103,106,109,96,96,97,103,102,105,110,109,88,93,97,100,100,107,115,114,90,93,97,98,102,105,109,113,82,83,92,95,97,99,107,114,63,73,86,85,92,91,98,102);
		wait for 10 ns;
		t_blur_matrix_int <= (103,98,101,102,98,100,108,112,107,105,105,111,109,112,118,123,108,112,114,125,121,118,117,131,108,115,121,127,133,129,126,131,113,121,125,133,141,141,138,134,114,117,121,126,142,145,141,140,112,117,118,118,130,137,137,141,105,110,113,117,125,124,136,140);
		wait for 10 ns;
		t_blur_matrix_int <= (113,115,120,121,117,119,122,123,127,134,140,135,128,126,126,128,139,139,145,145,137,131,125,129,142,148,145,140,142,134,137,135,138,143,138,137,144,141,141,134,144,138,142,137,145,151,148,133,146,146,142,140,140,142,139,128,139,145,134,133,135,133,131,122);
		wait for 10 ns;
		t_blur_matrix_int <= (126,118,103,112,110,73,14,43,124,117,114,115,110,30,18,46,124,118,116,121,81,10,20,34,125,117,124,116,47,17,29,35,119,116,125,103,20,17,37,29,117,122,121,75,16,20,38,27,114,120,108,62,15,19,34,27,113,114,103,64,18,23,36,37);
		wait for 10 ns;
		t_blur_matrix_int <= (27,21,19,21,21,29,27,30,24,15,20,25,24,27,26,38,22,20,23,25,23,30,36,33,18,22,24,24,29,33,37,29,22,28,30,23,30,29,38,35,31,32,31,29,31,29,35,39,33,36,35,32,31,33,36,45,37,37,36,36,34,31,43,42);
		wait for 10 ns;
		t_blur_matrix_int <= (32,34,25,26,20,21,20,68,30,39,23,29,19,23,24,76,44,28,22,27,24,23,26,83,37,19,36,33,17,23,31,79,32,19,42,25,23,25,36,86,23,18,32,23,22,24,35,83,21,29,24,27,24,24,43,86,29,38,23,28,25,28,46,81);
		wait for 10 ns;
		t_blur_matrix_int <= (51,48,54,54,41,34,33,58,53,44,54,55,47,40,45,53,55,48,62,49,44,38,45,56,57,50,63,57,38,39,46,50,62,50,68,54,40,48,47,42,60,53,70,48,43,56,47,45,61,47,67,45,40,54,47,48,64,59,64,53,46,59,55,51);
		wait for 10 ns;
		t_blur_matrix_int <= (36,18,26,44,132,147,126,138,38,21,30,33,131,152,134,142,40,26,30,32,131,153,134,143,36,37,25,36,133,148,135,144,35,46,22,26,136,152,135,138,38,47,34,27,132,157,135,142,33,51,25,28,135,149,134,143,45,55,32,34,136,145,131,136);
		wait for 10 ns;
		t_blur_matrix_int <= (124,123,138,133,138,138,137,135,120,127,137,138,138,141,141,138,117,134,134,143,139,139,137,139,116,131,133,144,139,140,135,139,121,130,134,143,139,141,138,131,120,128,137,139,139,140,138,135,124,129,130,133,137,136,135,134,120,116,117,122,124,126,127,127);
		wait for 10 ns;
		t_blur_matrix_int <= (135,134,137,135,136,133,135,135,136,134,138,134,134,132,132,135,137,135,137,134,133,134,132,133,134,137,135,133,132,134,131,136,131,133,133,132,132,132,131,132,130,130,134,132,134,134,133,129,129,135,133,131,133,133,132,131,129,134,128,135,131,133,131,129);
		wait for 10 ns;
		t_blur_matrix_int <= (135,134,130,131,129,130,128,126,135,136,131,134,129,131,126,128,138,136,130,131,132,129,125,127,135,134,134,134,133,130,128,124,133,135,129,131,129,130,123,125,134,130,133,132,133,129,126,124,134,133,132,130,126,125,125,124,128,131,130,129,127,124,125,121);
		wait for 10 ns;
		t_blur_matrix_int <= (126,124,125,122,120,114,107,102,127,124,124,120,118,113,105,104,124,122,122,122,119,113,107,101,126,123,123,120,117,115,109,103,123,122,122,118,115,113,108,104,123,121,119,121,118,113,109,99,121,119,119,119,114,109,105,98,121,123,117,118,118,110,104,98);
		wait for 10 ns;
		t_blur_matrix_int <= (98,102,151,192,210,213,214,214,97,100,158,193,208,215,214,214,95,105,162,196,210,214,214,214,96,113,172,201,214,216,214,213,95,118,180,205,214,217,215,212,98,126,184,208,217,219,214,210,99,137,190,209,219,219,211,208,101,152,195,211,217,214,214,208);
		wait for 10 ns;
		t_blur_matrix_int <= (210,209,208,211,211,211,210,211,211,211,209,210,210,208,207,208,211,208,208,208,206,205,207,206,210,209,207,205,207,205,206,207,207,205,206,205,206,206,209,209,205,205,205,205,208,208,208,209,205,204,206,207,208,210,211,210,204,205,207,207,207,208,208,208);
		wait for 10 ns;
		t_blur_matrix_int <= (208,207,203,203,202,203,204,204,208,205,205,204,206,208,205,207,206,206,206,207,205,205,209,203,211,207,208,207,206,204,202,203,209,209,207,205,203,200,201,199,209,209,205,203,202,197,197,199,208,206,202,201,198,199,199,195,205,205,200,200,198,196,194,190);
		wait for 10 ns;
		t_blur_matrix_int <= (203,205,202,204,204,205,204,204,204,206,203,203,202,203,202,200,201,202,200,201,201,199,196,199,202,200,200,200,198,199,198,195,198,197,198,199,197,198,196,192,196,195,195,195,192,187,180,170,195,189,185,180,169,157,134,103,187,175,155,133,102,69,46,28);
		wait for 10 ns;
		t_blur_matrix_int <= (16,19,23,22,21,18,15,26,23,17,23,24,17,17,20,19,20,22,24,21,20,15,16,15,28,32,29,29,18,15,16,17,30,34,35,33,26,20,20,16,43,42,40,37,29,24,26,21,78,66,53,43,37,29,27,22,107,98,82,67,53,46,36,29);
		wait for 10 ns;
		t_blur_matrix_int <= (20,28,48,68,70,73,91,102,17,30,45,66,64,64,84,101,16,28,45,59,60,57,72,96,15,28,40,50,48,49,79,100,13,26,32,47,47,46,75,99,18,24,34,40,36,43,66,87,22,30,35,36,28,33,52,78,27,35,25,28,19,26,40,66);
		wait for 10 ns;
		t_blur_matrix_int <= (118,128,136,144,151,150,152,152,112,127,135,144,151,152,150,151,112,125,134,143,150,153,149,153,111,125,133,147,151,152,152,152,108,122,133,142,149,150,149,151,103,116,130,143,148,148,150,146,96,115,131,141,150,149,146,147,87,111,129,141,146,147,151,146);
		wait for 10 ns;
		t_blur_matrix_int <= (157,157,157,152,146,131,112,91,153,156,159,152,140,132,109,83,154,154,153,151,139,129,107,81,149,151,153,152,142,123,103,81,150,155,157,149,139,122,106,105,149,150,154,145,136,126,127,172,149,146,154,147,142,140,179,140,148,150,151,159,176,155,127,90);
		wait for 10 ns;
		t_blur_matrix_int <= (65,38,25,46,102,93,57,85,61,32,55,129,176,76,85,116,55,66,153,189,75,35,82,98,86,158,190,72,78,37,101,76,171,177,67,48,38,32,90,42,145,51,36,56,34,60,121,21,68,34,36,48,41,126,86,16,64,39,43,75,114,109,36,16);
		wait for 10 ns;
		t_blur_matrix_int <= (24,20,44,74,44,47,34,36,19,20,31,56,46,29,39,34,24,14,24,61,53,30,36,38,32,31,17,58,56,42,38,39,18,17,20,55,66,44,30,41,19,17,13,41,67,42,31,38,15,18,11,31,59,46,18,35,17,19,16,20,35,59,40,59);
		wait for 10 ns;
		t_blur_matrix_int <= (38,38,44,34,22,25,29,14,32,46,25,28,23,26,23,15,35,42,24,30,21,22,19,14,50,27,30,49,23,22,24,19,41,32,30,68,34,32,29,23,39,30,30,69,58,34,27,25,27,24,27,71,77,40,42,37,12,18,22,48,82,54,49,36);
		wait for 10 ns;
		t_blur_matrix_int <= (67,141,117,95,39,52,54,42,52,138,127,128,74,76,63,36,47,123,108,137,106,54,56,38,62,118,101,103,128,78,56,46,51,107,109,89,120,125,69,38,38,61,105,114,82,109,119,55,35,23,55,119,96,65,108,102,62,13,20,99,113,96,55,41);
		wait for 10 ns;
		t_blur_matrix_int <= (67,94,104,69,95,123,83,109,54,103,119,74,59,99,83,110,32,72,118,66,53,111,111,61,24,38,69,64,91,141,112,62,18,34,87,100,119,141,80,66,42,57,79,120,146,107,48,73,111,116,119,147,133,51,62,60,65,76,107,142,70,54,70,79);
		wait for 10 ns;
		t_blur_matrix_int <= (116,141,134,104,120,104,110,48,131,146,122,112,135,153,144,101,123,140,125,83,49,78,134,145,81,136,146,119,64,32,54,148,82,101,127,84,104,71,32,94,69,70,101,112,67,63,56,73,91,73,78,113,87,46,103,115,63,98,93,89,90,80,102,139);
		wait for 10 ns;
		t_blur_matrix_int <= (25,22,25,27,27,28,29,27,40,30,28,30,28,29,30,28,96,47,20,17,22,23,28,22,162,131,47,21,22,23,23,25,148,148,131,48,26,28,27,30,135,106,140,130,35,20,24,31,147,101,53,153,104,30,20,27,149,83,54,66,147,56,19,25);
		wait for 10 ns;
		t_blur_matrix_int <= (29,38,46,38,19,20,33,45,32,50,48,41,24,20,29,45,28,47,51,38,18,15,31,36,28,44,55,33,18,15,42,38,35,45,59,29,22,23,45,46,41,43,56,31,22,21,36,46,26,40,48,23,18,21,43,49,28,40,53,22,23,23,44,50);
		wait for 10 ns;
		t_blur_matrix_int <= (26,24,22,28,30,22,22,24,24,27,24,24,32,23,23,27,24,24,24,23,28,24,22,27,22,22,21,22,29,27,22,25,23,23,28,22,28,29,22,20,30,28,30,23,20,25,33,27,24,26,29,24,23,23,30,27,20,24,23,19,26,19,31,26);
		wait for 10 ns;
		t_blur_matrix_int <= (16,21,27,27,34,32,30,39,23,21,27,26,33,38,33,34,22,21,26,24,30,36,34,29,23,19,26,22,32,31,34,26,23,21,24,24,29,31,35,28,21,29,28,29,24,26,36,36,23,26,25,23,26,22,33,34,24,22,25,19,23,31,36,38);
		wait for 10 ns;
		t_blur_matrix_int <= (37,39,29,32,43,43,43,33,37,37,32,26,31,39,55,45,33,31,32,25,25,38,44,45,37,30,25,21,21,36,43,51,29,34,29,22,23,26,46,50,27,31,28,30,22,30,50,55,31,30,31,28,24,24,41,56,31,33,30,31,24,19,40,53);
		wait for 10 ns;
		t_blur_matrix_int <= (27,27,23,30,27,34,32,34,33,30,35,47,46,53,53,61,48,50,61,77,79,81,91,96,53,65,76,79,89,93,96,94,57,69,79,86,95,96,94,88,57,74,84,90,93,95,89,91,62,76,79,88,87,90,91,90,60,78,88,88,85,90,89,92);
		wait for 10 ns;
		t_blur_matrix_int <= (39,47,59,64,77,83,89,91,71,73,76,76,80,85,92,88,98,101,111,111,106,104,109,112,95,99,108,105,104,105,107,111,95,96,97,101,100,104,104,106,93,95,102,98,100,103,107,105,89,89,94,98,100,106,103,104,91,90,91,95,106,104,101,102);
		wait for 10 ns;
		t_blur_matrix_int <= (100,106,109,119,120,116,125,136,95,99,99,118,116,124,122,128,110,117,117,134,130,137,130,133,106,108,116,122,126,129,125,122,109,112,117,118,120,124,118,121,103,109,112,117,118,116,113,112,106,107,112,114,113,107,113,107,103,106,108,109,105,110,107,111);
		wait for 10 ns;
		t_blur_matrix_int <= (137,138,131,123,120,123,123,112,140,137,130,126,125,123,113,104,136,143,142,147,149,148,147,149,128,127,130,130,132,136,147,155,116,118,119,121,129,135,148,159,115,113,113,117,127,138,154,158,112,113,113,124,127,148,149,161,112,111,115,123,133,145,151,166);
		wait for 10 ns;
		t_blur_matrix_int <= (112,107,94,48,23,23,27,31,104,109,85,51,29,30,29,34,154,157,142,97,64,46,34,39,165,178,183,183,172,143,92,56,169,180,183,185,188,189,188,162,168,180,186,186,188,189,192,194,173,179,186,186,189,191,188,192,174,178,184,184,187,187,191,191);
		wait for 10 ns;
		t_blur_matrix_int <= (33,30,35,35,32,29,43,32,39,40,31,37,33,28,43,36,40,34,35,32,33,30,35,33,34,35,31,35,27,26,28,32,107,63,43,39,31,27,26,32,191,169,116,69,42,33,30,30,191,192,192,177,123,62,31,24,192,189,192,196,197,177,118,53);
		wait for 10 ns;
		t_blur_matrix_int <= (28,30,28,22,29,36,46,79,33,25,27,26,23,36,44,78,32,24,28,27,25,37,41,76,26,21,25,33,22,39,40,74,23,21,22,26,27,45,48,71,32,25,27,27,28,40,62,72,23,15,19,13,23,32,61,56,23,15,15,11,18,31,48,58);
		wait for 10 ns;
		t_blur_matrix_int <= (66,62,61,56,47,61,58,53,64,60,67,61,52,52,56,53,73,55,69,57,49,57,57,47,70,55,70,57,51,52,59,56,74,50,59,66,51,48,57,54,79,53,62,59,47,51,61,52,79,47,57,55,46,46,59,51,80,39,58,56,50,43,57,42);
		wait for 10 ns;
		t_blur_matrix_int <= (38,55,32,40,141,143,135,129,37,47,42,43,142,142,137,121,41,43,43,51,150,134,137,109,43,43,38,58,148,127,132,101,48,48,42,63,152,128,128,98,42,55,44,71,158,126,119,98,38,51,35,80,154,126,115,102,41,36,35,87,146,124,115,107);
		wait for 10 ns;
		t_blur_matrix_int <= (112,104,102,107,114,118,116,122,102,96,89,93,99,105,109,108,88,97,83,85,89,96,97,98,80,93,88,79,83,83,89,90,90,92,99,89,85,88,82,91,98,109,104,106,92,97,89,88,108,113,108,112,109,101,102,97,115,115,113,114,117,107,105,105);
		wait for 10 ns;
		t_blur_matrix_int <= (127,124,128,133,130,132,135,132,116,113,116,119,125,125,123,126,102,109,104,110,115,116,118,118,93,96,90,97,98,102,106,108,87,85,89,90,89,91,92,97,86,85,83,83,80,83,84,84,92,91,86,84,79,80,78,79,101,100,93,88,87,82,77,75);
		wait for 10 ns;
		t_blur_matrix_int <= (134,130,129,128,128,127,125,124,130,132,129,127,128,127,125,122,125,129,129,128,126,125,124,121,112,115,120,121,119,120,121,121,101,103,106,109,111,113,116,117,87,83,94,94,94,99,97,105,76,75,81,85,88,90,88,87,74,73,74,68,72,80,74,75);
		wait for 10 ns;
		t_blur_matrix_int <= (125,121,117,119,115,109,99,96,121,118,115,116,108,106,98,95,120,120,115,112,109,104,96,96,120,120,114,112,104,102,97,101,115,117,114,109,108,102,96,99,106,108,106,105,101,101,95,100,91,91,92,92,93,89,84,96,77,76,83,89,81,71,68,85);
		wait for 10 ns;
		t_blur_matrix_int <= (111,168,197,213,215,213,210,207,119,178,201,212,216,210,207,205,138,188,207,211,213,207,204,202,151,191,208,213,209,201,199,202,157,196,207,209,204,198,199,199,160,194,205,208,202,195,196,199,160,192,204,202,197,195,196,199,149,186,200,200,197,193,197,199);
		wait for 10 ns;
		t_blur_matrix_int <= (204,206,204,206,208,206,206,202,204,205,205,204,203,205,202,203,203,203,205,200,202,203,200,199,202,203,205,200,201,199,199,196,199,203,201,202,199,199,195,191,200,202,200,201,202,201,192,184,201,202,203,201,203,200,192,179,199,199,200,202,199,198,190,171);
		wait for 10 ns;
		t_blur_matrix_int <= (203,200,200,199,193,189,180,170,201,200,194,187,183,168,146,118,199,192,183,172,157,132,89,47,194,187,173,155,137,100,56,21,187,180,166,148,112,68,30,21,174,167,149,122,75,30,15,15,167,145,101,61,30,15,14,22,150,101,43,19,21,22,28,37);
		wait for 10 ns;
		t_blur_matrix_int <= (154,127,85,47,23,20,21,18,76,45,24,21,12,16,19,19,24,17,17,17,16,21,26,28,17,19,19,23,19,34,46,42,15,15,19,31,41,48,52,47,20,31,32,42,48,55,54,51,30,32,41,49,54,56,53,63,37,41,42,55,53,52,58,59);
		wait for 10 ns;
		t_blur_matrix_int <= (113,112,107,95,72,61,52,39,123,116,116,113,97,83,64,54,122,117,126,121,114,102,87,76,119,116,124,130,132,122,108,92,110,118,127,135,138,130,125,109,108,116,125,131,140,137,136,122,108,105,114,129,139,140,139,131,74,81,108,120,130,138,147,140);
		wait for 10 ns;
		t_blur_matrix_int <= (34,44,31,25,21,23,37,62,49,52,39,30,23,21,40,62,64,63,50,34,19,15,40,61,75,67,56,38,19,19,31,60,95,79,59,39,24,13,31,61,110,95,71,46,32,15,36,59,119,116,87,60,31,15,34,55,138,129,102,65,31,15,33,64);
		wait for 10 ns;
		t_blur_matrix_int <= (84,109,127,139,146,145,148,150,84,110,130,139,143,146,144,149,81,110,130,139,144,145,147,147,87,110,126,140,143,149,147,147,88,110,129,145,150,153,151,150,84,109,132,141,153,152,154,152,86,111,132,141,153,156,153,152,87,110,128,144,155,154,155,156);
		wait for 10 ns;
		t_blur_matrix_int <= (150,148,159,167,154,135,116,93,147,144,153,149,146,134,115,92,147,150,150,150,141,132,114,89,150,151,153,148,143,127,109,95,148,151,157,151,141,129,106,123,152,152,156,151,141,127,109,147,150,152,157,149,140,126,113,156,156,154,159,154,143,131,111,128);
		wait for 10 ns;
		t_blur_matrix_int <= (66,45,76,96,169,40,17,16,67,68,103,119,138,21,22,18,100,117,94,122,72,21,16,22,134,164,66,93,46,19,21,22,198,147,62,64,49,34,20,16,206,111,83,59,26,29,27,22,203,88,110,120,12,16,13,24,180,65,71,101,15,16,22,20);
		wait for 10 ns;
		t_blur_matrix_int <= (16,17,15,20,18,46,79,73,18,20,20,16,26,38,82,72,15,15,14,14,60,85,89,68,21,14,12,9,22,73,99,111,17,14,18,18,22,41,33,37,25,24,24,22,36,54,22,17,32,33,30,36,39,52,33,20,26,27,20,28,49,36,43,29);
		wait for 10 ns;
		t_blur_matrix_int <= (6,15,23,37,96,69,48,56,10,13,17,38,111,68,49,82,22,14,26,83,118,47,54,71,98,87,108,106,55,45,45,45,59,87,76,48,45,55,33,39,40,52,40,38,33,25,35,53,47,54,36,28,36,40,38,32,24,34,18,24,58,62,39,31);
		wait for 10 ns;
		t_blur_matrix_int <= (67,12,10,34,98,119,102,73,64,25,15,22,52,91,97,118,37,28,16,44,76,51,33,74,58,17,43,96,65,33,40,94,47,65,101,83,23,18,50,121,67,66,58,34,11,19,92,123,25,21,30,33,25,27,86,103,19,18,19,54,33,18,32,66);
		wait for 10 ns;
		t_blur_matrix_int <= (66,57,87,112,34,85,84,76,83,82,123,84,46,44,98,91,93,121,75,39,49,54,48,102,104,58,53,35,50,62,58,63,45,33,45,34,34,62,78,59,27,36,39,54,42,42,75,80,49,24,40,58,53,48,55,89,86,37,29,43,41,54,46,66);
		wait for 10 ns;
		t_blur_matrix_int <= (84,76,102,102,93,88,97,102,91,89,64,135,105,104,117,97,102,95,72,111,140,104,115,88,96,105,101,133,126,126,115,117,82,97,109,118,120,121,127,141,65,68,91,117,117,113,147,129,74,64,75,111,128,115,125,98,92,70,61,108,126,115,115,95);
		wait for 10 ns;
		t_blur_matrix_int <= (146,67,58,47,68,124,34,27,104,134,45,24,82,118,87,24,76,111,122,26,31,76,134,44,38,28,102,95,25,46,109,108,68,12,66,161,71,26,63,155,123,26,20,127,162,42,69,116,119,86,45,86,155,114,68,64,105,120,77,89,82,131,57,29);
		wait for 10 ns;
		t_blur_matrix_int <= (23,38,47,23,20,14,42,44,27,40,40,24,17,14,52,44,28,37,28,25,20,20,51,46,25,34,33,30,26,25,52,46,39,28,30,21,20,22,48,43,80,22,19,19,22,21,44,44,141,32,26,23,30,30,50,45,163,52,24,22,23,21,52,39);
		wait for 10 ns;
		t_blur_matrix_int <= (20,23,23,19,23,18,28,31,27,26,33,22,25,18,32,29,24,29,28,27,28,24,26,31,29,30,30,26,25,23,31,31,29,28,27,31,29,25,29,31,25,29,25,27,31,28,26,31,32,35,33,35,35,32,34,36,37,37,26,23,28,19,25,34);
		wait for 10 ns;
		t_blur_matrix_int <= (29,26,23,20,27,32,28,35,37,34,28,23,27,26,28,32,38,43,28,29,27,28,30,33,36,36,34,28,25,24,35,37,40,38,28,28,27,24,39,33,39,39,26,25,31,30,46,42,39,46,33,34,35,34,53,48,35,43,30,30,25,23,36,40);
		wait for 10 ns;
		t_blur_matrix_int <= (33,47,32,27,25,21,32,48,36,43,39,31,27,24,33,52,33,45,51,34,29,26,31,54,37,35,54,36,27,29,28,57,38,44,58,53,31,20,23,56,32,48,63,66,34,20,19,47,34,54,70,72,48,27,19,46,36,54,76,76,55,21,16,38);
		wait for 10 ns;
		t_blur_matrix_int <= (62,71,80,82,87,89,88,86,67,72,78,78,81,89,88,91,66,70,84,80,82,85,87,91,63,76,80,82,83,83,92,92,57,80,80,80,88,93,89,90,53,83,81,79,85,96,85,79,56,89,87,84,82,87,78,87,55,89,88,79,77,83,95,93);
		wait for 10 ns;
		t_blur_matrix_int <= (91,90,95,93,103,103,99,99,93,95,94,94,97,102,101,107,90,95,90,96,100,104,105,110,90,90,97,97,100,105,110,112,83,89,103,104,102,99,104,110,87,98,102,108,103,99,101,105,102,97,98,106,101,103,105,109,97,98,103,104,104,108,106,105);
		wait for 10 ns;
		t_blur_matrix_int <= (103,106,107,104,111,106,107,111,104,110,107,106,109,105,109,114,107,108,107,104,106,100,109,114,108,107,110,98,102,101,109,113,108,108,107,102,103,106,107,115,104,108,106,107,105,110,113,118,111,104,104,105,107,112,118,119,111,104,110,107,108,114,118,120);
		wait for 10 ns;
		t_blur_matrix_int <= (113,117,119,128,136,150,159,171,112,118,125,132,140,150,158,166,115,120,128,134,147,154,160,165,117,126,131,138,140,148,151,163,122,128,133,138,142,144,149,160,124,128,133,137,139,144,149,157,126,131,138,135,143,145,147,144,124,131,137,134,138,140,145,150);
		wait for 10 ns;
		t_blur_matrix_int <= (175,177,179,184,181,186,187,189,173,175,177,175,179,183,183,185,171,177,176,174,178,182,183,181,168,173,171,174,177,178,178,179,162,168,166,170,177,174,177,179,158,161,163,166,171,172,175,178,155,156,164,159,163,175,173,173,156,154,157,157,165,162,166,167);
		wait for 10 ns;
		t_blur_matrix_int <= (191,193,191,194,194,198,199,169,189,191,189,192,192,198,201,201,187,190,191,193,194,196,198,199,185,186,190,192,191,195,197,198,183,186,184,191,192,195,197,198,182,180,183,187,189,194,194,197,180,178,183,186,190,192,196,196,174,181,183,185,188,191,194,194);
		wait for 10 ns;
		t_blur_matrix_int <= (86,35,18,12,18,37,45,60,191,126,44,17,17,33,29,58,202,201,154,58,25,28,22,49,200,203,204,166,64,26,17,36,201,202,203,207,172,68,19,31,198,201,202,206,207,170,58,31,197,201,200,208,208,208,158,44,197,201,201,204,207,210,210,135);
		wait for 10 ns;
		t_blur_matrix_int <= (79,44,55,52,46,39,52,43,76,36,48,52,42,43,48,39,74,40,50,53,40,48,56,39,65,34,40,43,34,40,52,41,58,29,33,37,31,44,47,41,52,34,35,34,39,54,49,44,32,29,21,27,32,45,33,47,30,21,13,18,29,45,34,36);
		wait for 10 ns;
		t_blur_matrix_int <= (43,39,36,94,142,122,118,117,47,32,35,109,140,120,111,124,44,25,37,122,133,120,113,126,40,21,35,132,127,116,116,134,35,16,33,132,129,117,116,130,41,20,47,140,124,119,119,128,44,17,51,148,117,119,118,126,33,18,64,147,113,116,124,129);
		wait for 10 ns;
		t_blur_matrix_int <= (123,118,117,117,121,114,112,110,125,126,120,121,120,120,114,114,128,124,126,125,121,119,118,116,128,125,124,125,124,123,120,121,127,129,123,127,123,122,121,124,130,131,125,126,125,124,129,120,130,130,127,128,125,118,124,123,131,129,127,125,125,121,123,120);
		wait for 10 ns;
		t_blur_matrix_int <= (108,105,103,102,98,89,86,85,114,114,109,109,106,103,97,93,115,116,116,113,110,105,104,98,119,119,116,113,117,111,110,107,121,125,119,114,115,114,113,108,124,121,119,121,119,116,118,115,122,123,120,118,119,116,117,114,122,123,119,121,119,119,116,113);
		wait for 10 ns;
		t_blur_matrix_int <= (80,75,71,70,68,73,71,65,89,87,78,76,71,73,64,64,101,93,91,82,83,83,73,64,105,98,95,97,89,87,82,71,106,103,103,99,96,95,95,82,110,107,112,106,104,105,97,92,113,110,108,108,105,106,100,99,114,113,109,110,107,109,102,103);
		wait for 10 ns;
		t_blur_matrix_int <= (72,75,86,89,80,63,48,68,70,82,99,96,87,66,48,61,78,87,107,102,83,67,43,70,79,91,105,106,89,66,50,93,88,99,107,106,86,69,60,119,95,102,103,106,91,78,78,140,95,101,105,105,100,84,95,158,102,103,113,108,99,91,117,176);
		wait for 10 ns;
		t_blur_matrix_int <= (139,186,199,199,195,194,200,202,141,189,200,200,197,197,202,204,150,189,200,203,199,200,205,206,162,195,203,202,203,204,205,206,180,196,204,206,206,204,206,206,186,201,206,204,205,206,205,205,193,203,206,207,205,206,206,205,196,207,205,207,206,208,206,204);
		wait for 10 ns;
		t_blur_matrix_int <= (202,199,199,199,193,187,177,150,201,199,199,197,184,166,146,103,203,201,199,194,170,132,85,36,203,200,197,191,154,92,35,25,201,196,192,176,128,67,19,16,200,193,182,160,111,41,14,23,200,189,170,137,88,29,24,39,198,180,155,112,68,32,39,57);
		wait for 10 ns;
		t_blur_matrix_int <= (116,53,15,19,29,41,43,43,55,25,18,37,44,50,51,47,16,18,35,47,54,49,48,51,16,33,58,58,53,48,47,49,33,58,63,60,57,55,50,57,48,58,61,63,57,53,54,66,62,61,60,64,65,58,60,77,66,62,56,61,61,63,72,80);
		wait for 10 ns;
		t_blur_matrix_int <= (42,48,51,55,54,56,56,54,53,52,55,60,60,54,61,56,58,59,63,62,64,56,50,55,59,63,67,68,61,55,50,56,68,70,73,67,62,58,53,63,73,75,72,66,60,61,59,69,83,85,75,66,61,51,65,64,83,76,71,66,61,63,70,74);
		wait for 10 ns;
		t_blur_matrix_int <= (41,58,92,113,125,138,154,152,20,39,74,102,119,143,154,153,12,24,57,88,114,146,151,157,9,17,29,67,106,142,158,162,7,9,22,52,109,140,158,159,12,13,21,46,96,139,160,163,10,18,21,38,88,136,153,163,7,10,22,44,86,129,149,160);
		wait for 10 ns;
		t_blur_matrix_int <= (149,132,113,79,32,15,29,58,153,139,119,92,47,12,29,56,157,141,123,101,49,11,24,56,162,148,133,112,52,14,17,49,159,150,135,111,56,9,11,43,161,157,144,113,40,12,15,46,164,156,142,105,43,13,13,50,162,156,137,105,46,7,10,42);
		wait for 10 ns;
		t_blur_matrix_int <= (86,115,132,144,156,156,156,154,88,112,130,143,158,154,154,156,89,117,131,147,152,157,159,158,86,116,130,145,155,153,153,155,91,113,131,143,152,159,159,153,87,116,133,140,158,160,158,158,86,115,129,144,156,161,161,157,87,112,132,146,158,156,158,157);
		wait for 10 ns;
		t_blur_matrix_int <= (154,159,161,152,143,129,113,135,156,160,157,153,144,126,118,142,154,157,160,152,143,132,115,116,158,160,157,153,143,133,119,99,153,157,160,157,146,135,120,99,156,160,158,154,148,138,123,99,158,160,159,157,150,138,124,103,156,160,162,159,151,136,120,102);
		wait for 10 ns;
		t_blur_matrix_int <= (126,88,47,32,16,16,24,16,154,94,50,34,19,18,21,17,158,88,64,55,15,13,22,15,90,146,74,47,12,18,26,18,80,145,50,26,19,24,19,18,75,86,113,19,19,26,23,17,101,94,104,23,29,22,20,25,148,100,63,24,30,16,19,34);
		wait for 10 ns;
		t_blur_matrix_int <= (18,26,20,30,51,24,35,30,16,26,22,60,37,23,34,27,24,21,29,70,24,27,22,42,19,27,50,40,23,19,26,31,33,33,37,28,20,22,28,26,23,38,31,26,23,24,26,25,38,34,26,29,24,23,27,28,37,25,19,26,15,15,26,26);
		wait for 10 ns;
		t_blur_matrix_int <= (22,22,16,25,73,75,33,44,27,18,17,37,84,69,19,60,27,23,18,40,95,70,20,49,23,25,19,40,102,75,21,43,17,19,22,44,108,65,16,38,23,21,19,60,126,57,15,28,25,26,22,86,126,56,13,16,20,19,36,115,116,49,15,15);
		wait for 10 ns;
		t_blur_matrix_int <= (25,20,18,60,55,17,20,49,35,16,13,40,84,29,17,40,34,13,12,20,73,51,19,29,43,20,14,13,30,65,44,23,56,23,13,12,16,27,69,58,61,23,12,21,29,24,37,61,56,41,13,29,30,17,38,27,42,38,12,40,34,23,45,27);
		wait for 10 ns;
		t_blur_matrix_int <= (84,71,27,36,50,51,44,52,62,59,67,33,46,57,54,51,72,36,63,65,36,75,71,56,68,34,42,76,62,63,81,87,62,46,24,49,65,59,81,92,68,58,26,53,44,71,71,91,26,37,20,58,38,72,68,81,14,29,28,46,51,55,78,81);
		wait for 10 ns;
		t_blur_matrix_int <= (81,89,61,107,128,110,111,123,49,91,67,104,90,91,98,128,40,58,72,104,63,94,106,100,76,50,61,91,62,110,114,88,93,73,48,68,58,101,121,131,83,74,57,67,53,85,135,141,73,69,52,65,56,85,124,138,94,75,62,52,50,90,126,120);
		wait for 10 ns;
		t_blur_matrix_int <= (110,134,68,98,37,119,133,25,120,160,120,91,18,42,167,58,123,157,144,74,17,14,81,94,122,155,135,82,34,9,37,122,115,144,100,26,41,17,37,142,125,140,131,30,21,56,23,133,118,130,141,61,20,27,21,126,93,141,116,94,30,20,16,119);
		wait for 10 ns;
		t_blur_matrix_int <= (148,100,14,14,19,15,50,36,128,142,16,12,16,17,44,35,116,171,17,10,13,13,41,38,121,194,24,21,16,13,41,37,146,195,32,17,14,15,46,34,167,182,17,12,12,12,48,29,180,148,18,14,20,21,55,38,176,86,27,9,12,23,58,32);
		wait for 10 ns;
		t_blur_matrix_int <= (28,33,23,22,25,20,24,26,30,38,24,27,24,24,26,27,29,39,22,23,23,18,21,29,30,47,23,23,20,19,27,25,32,50,25,25,23,24,25,32,37,64,22,23,22,21,24,25,35,65,28,29,27,31,22,28,39,53,20,32,25,21,24,24);
		wait for 10 ns;
		t_blur_matrix_int <= (37,46,25,23,21,16,35,41,36,36,34,29,27,16,34,40,51,42,27,30,39,17,28,29,39,47,26,30,28,19,30,28,41,34,21,22,26,17,25,27,38,34,23,23,34,29,26,41,40,30,18,18,23,23,28,49,41,40,26,18,20,29,26,57);
		wait for 10 ns;
		t_blur_matrix_int <= (36,62,80,83,70,23,16,33,34,63,85,81,69,32,15,35,36,67,83,84,72,38,9,27,50,76,81,82,69,33,11,24,58,66,73,83,63,40,17,23,64,78,73,62,68,48,16,25,69,72,63,71,79,47,17,26,61,63,70,89,83,54,17,26);
		wait for 10 ns;
		t_blur_matrix_int <= (56,81,84,70,79,98,102,92,54,75,71,76,91,98,99,93,48,72,85,83,88,97,100,98,52,75,80,82,92,98,94,96,58,69,83,81,92,94,88,94,59,71,84,86,92,95,89,90,62,67,80,90,98,94,92,92,65,72,82,92,95,92,92,96);
		wait for 10 ns;
		t_blur_matrix_int <= (92,100,104,103,104,104,108,103,94,99,101,102,106,107,107,102,98,91,100,100,102,108,107,109,97,99,98,99,103,105,109,105,101,99,95,96,102,101,107,107,96,100,100,102,104,102,107,105,97,103,103,104,104,102,102,104,105,101,100,103,102,103,98,101);
		wait for 10 ns;
		t_blur_matrix_int <= (102,105,103,109,113,109,116,120,105,104,105,110,108,113,111,120,109,108,106,107,110,108,117,119,106,108,109,109,112,113,114,118,109,106,107,108,116,117,120,119,105,108,107,110,115,117,115,113,105,107,109,111,106,113,116,112,103,103,105,104,110,115,113,113);
		wait for 10 ns;
		t_blur_matrix_int <= (121,124,135,135,133,137,143,145,121,122,125,136,134,137,141,141,123,124,130,132,135,137,137,142,117,120,125,128,135,133,142,140,117,122,126,126,131,134,137,138,120,118,122,129,129,132,135,136,115,122,126,128,127,131,131,133,115,119,123,126,125,130,130,138);
		wait for 10 ns;
		t_blur_matrix_int <= (153,158,154,156,157,166,166,167,147,154,154,157,163,160,165,173,148,148,151,153,160,160,165,169,142,145,152,155,159,159,168,163,144,148,150,153,155,161,163,163,139,146,152,152,155,160,158,169,143,143,149,149,156,154,161,170,141,142,147,151,150,156,161,162);
		wait for 10 ns;
		t_blur_matrix_int <= (173,180,181,183,187,189,193,195,172,177,177,181,183,186,191,192,172,176,177,182,184,188,189,191,172,178,178,181,184,187,190,194,169,174,174,180,184,185,191,190,169,175,174,177,186,187,188,194,170,169,173,177,181,187,190,193,167,173,173,179,181,183,187,190);
		wait for 10 ns;
		t_blur_matrix_int <= (197,200,200,205,207,209,210,204,195,197,198,204,204,209,211,215,192,197,197,202,203,207,211,216,195,196,197,202,204,205,210,214,194,197,200,201,201,206,209,211,196,198,199,205,202,204,207,211,195,199,196,203,202,203,208,210,194,196,196,201,204,204,205,207);
		wait for 10 ns;
		t_blur_matrix_int <= (100,29,17,18,23,38,23,37,185,60,20,18,22,30,18,32,214,145,19,13,21,49,15,33,215,201,69,20,14,22,14,24,213,216,149,17,14,19,11,15,213,215,201,59,12,16,9,13,212,213,215,133,10,9,7,10,211,215,216,192,31,17,8,9);
		wait for 10 ns;
		t_blur_matrix_int <= (22,14,73,147,114,116,126,127,24,18,92,135,107,119,119,128,16,18,106,129,109,119,125,130,10,19,113,127,107,116,131,129,9,26,120,137,109,119,132,129,6,31,128,132,109,124,132,131,5,46,121,131,113,125,128,130,6,62,121,123,121,127,130,129);
		wait for 10 ns;
		t_blur_matrix_int <= (128,127,126,128,126,123,125,120,126,127,130,124,124,124,127,126,128,126,124,125,123,127,128,122,125,128,125,124,121,121,126,120,125,123,124,127,124,123,125,123,129,128,125,127,122,125,124,124,132,133,124,125,129,126,122,123,127,130,126,128,124,125,121,120);
		wait for 10 ns;
		t_blur_matrix_int <= (120,123,120,124,119,121,117,116,124,122,123,123,120,120,119,117,120,124,119,119,120,118,119,117,120,119,120,118,119,116,118,118,119,122,119,121,116,115,115,119,121,119,119,118,114,114,114,114,123,124,117,120,117,115,115,115,123,119,120,115,110,111,112,112);
		wait for 10 ns;
		t_blur_matrix_int <= (114,113,114,109,108,106,105,106,113,119,114,110,106,105,111,103,116,117,112,112,108,111,109,102,115,116,114,110,112,106,102,101,115,113,115,109,106,103,103,95,115,112,113,107,101,104,97,97,115,110,110,107,103,102,98,111,113,110,108,103,100,100,98,128);
		wait for 10 ns;
		t_blur_matrix_int <= (104,108,114,113,104,94,132,185,106,112,112,114,112,106,146,189,101,108,110,117,117,118,163,192,97,104,123,137,149,160,177,195,102,120,138,157,170,179,192,201,115,141,161,178,183,188,198,203,142,166,181,187,189,193,199,209,173,189,197,195,190,193,200,209);
		wait for 10 ns;
		t_blur_matrix_int <= (201,208,208,205,208,205,205,202,206,212,208,206,208,206,207,200,207,211,207,206,208,204,201,200,207,209,207,209,207,204,203,198,208,210,209,207,206,204,198,191,210,211,208,210,205,200,197,179,211,210,210,208,205,199,189,162,213,210,210,209,205,196,178,138);
		wait for 10 ns;
		t_blur_matrix_int <= (196,173,129,87,48,39,51,65,191,162,110,61,44,45,59,67,187,148,85,45,45,54,61,63,178,125,67,46,53,59,62,57,158,104,57,54,56,65,64,56,137,76,58,59,63,65,61,65,105,64,56,62,62,61,65,69,87,58,60,61,59,57,68,73);
		wait for 10 ns;
		t_blur_matrix_int <= (66,58,61,63,65,69,79,81,62,62,68,66,70,79,85,86,57,69,70,67,73,84,83,73,64,70,75,78,82,81,70,66,67,70,75,80,82,79,66,62,70,72,76,83,80,74,67,61,75,76,81,85,76,67,62,59,77,82,85,85,71,62,63,57);
		wait for 10 ns;
		t_blur_matrix_int <= (82,76,68,63,58,64,72,75,75,63,63,64,65,77,74,76,66,59,62,65,72,72,77,74,57,56,60,74,73,74,71,76,55,58,63,73,74,76,75,74,62,63,67,75,73,70,75,78,62,67,71,77,72,67,77,80,64,74,73,72,72,72,83,81);
		wait for 10 ns;
		t_blur_matrix_int <= (7,7,9,30,82,131,143,158,5,8,8,24,74,122,146,158,9,8,8,19,65,117,147,161,5,8,9,25,66,116,146,162,6,8,7,19,68,119,143,157,8,6,8,15,63,114,141,157,7,6,9,17,57,106,145,158,9,7,9,16,49,100,141,153);
		wait for 10 ns;
		t_blur_matrix_int <= (162,159,141,110,48,7,14,40,162,160,143,114,48,9,11,37,163,159,144,115,57,8,11,34,168,161,143,120,66,11,10,34,165,159,144,120,72,16,11,35,164,160,149,121,86,20,13,32,164,161,149,126,84,15,11,35,165,162,155,133,81,21,15,33);
		wait for 10 ns;
		t_blur_matrix_int <= (83,113,131,144,155,162,158,160,86,113,134,148,157,159,159,159,85,111,133,146,159,161,158,157,81,111,129,149,155,158,158,155,79,113,132,146,160,155,156,157,77,109,130,146,154,156,151,151,74,109,130,146,155,157,156,155,78,107,133,146,153,154,158,159);
		wait for 10 ns;
		t_blur_matrix_int <= (158,159,163,159,151,137,122,100,159,162,165,154,145,138,119,105,162,162,163,160,150,137,124,103,159,160,161,159,152,136,124,105,158,157,157,155,145,135,125,112,152,148,150,154,145,133,124,106,154,153,160,155,146,132,120,108,159,157,161,156,149,140,122,117);
		wait for 10 ns;
		t_blur_matrix_int <= (142,94,57,21,28,19,27,41,125,71,18,21,29,27,33,29,113,70,22,25,34,36,29,13,98,67,28,37,37,25,21,19,90,75,39,37,33,18,21,21,102,107,39,24,29,19,22,24,114,98,38,39,18,19,21,21,109,70,33,29,27,23,19,32);
		wait for 10 ns;
		t_blur_matrix_int <= (27,22,23,20,22,17,30,13,20,16,17,18,19,22,21,11,21,18,20,17,21,22,13,17,22,23,23,16,21,20,19,28,25,19,21,20,23,22,41,49,16,21,30,24,22,52,69,26,20,19,28,26,20,41,35,22,20,22,27,19,22,23,22,32);
		wait for 10 ns;
		t_blur_matrix_int <= (12,19,72,112,106,46,22,24,10,41,121,102,100,48,18,16,37,94,90,68,74,28,18,18,99,70,28,78,65,46,24,18,46,19,26,97,60,49,26,22,24,21,30,66,59,61,21,28,28,27,28,67,61,51,26,24,35,24,25,55,54,41,28,25);
		wait for 10 ns;
		t_blur_matrix_int <= (27,36,16,51,30,28,28,36,19,31,22,44,27,31,15,24,21,25,41,44,17,30,12,12,24,33,52,38,17,31,14,15,20,32,55,35,18,21,21,17,17,41,33,39,23,21,23,20,36,37,21,37,24,27,24,26,41,27,20,35,34,24,20,17);
		wait for 10 ns;
		t_blur_matrix_int <= (20,29,22,27,50,48,62,80,20,33,24,22,42,41,51,64,23,41,32,14,47,37,37,36,19,40,36,8,40,45,31,57,23,38,39,11,40,64,29,26,24,47,22,25,43,65,36,23,19,42,29,29,65,64,28,23,18,37,32,23,80,55,17,44);
		wait for 10 ns;
		t_blur_matrix_int <= (99,72,54,52,37,83,144,109,112,89,31,33,38,88,137,122,100,102,40,47,68,100,122,123,99,90,92,75,85,102,120,123,46,51,93,108,114,106,114,135,22,30,57,105,128,111,100,125,11,21,53,101,132,101,114,112,15,32,52,90,107,73,129,79);
		wait for 10 ns;
		t_blur_matrix_int <= (105,143,109,124,96,41,32,140,131,144,65,77,124,72,107,164,137,145,121,67,113,53,135,150,122,75,119,121,129,140,174,123,105,54,75,109,117,145,149,127,109,85,61,58,81,115,97,142,112,70,72,10,11,47,48,28,98,107,89,48,12,31,70,16);
		wait for 10 ns;
		t_blur_matrix_int <= (141,59,115,14,13,26,55,36,119,125,176,28,14,29,44,31,108,113,94,18,19,33,39,23,29,18,14,37,33,40,30,25,88,37,38,67,21,43,28,29,151,119,118,81,62,70,37,32,35,63,70,82,112,107,91,115,20,48,10,18,45,48,37,99);
		wait for 10 ns;
		t_blur_matrix_int <= (44,41,24,30,25,25,19,28,39,33,32,26,34,29,23,23,31,34,38,26,33,33,25,34,34,29,35,21,32,29,23,35,38,28,37,32,35,28,24,34,30,32,48,57,30,25,30,31,94,89,61,31,32,22,22,30,91,74,80,46,32,25,33,28);
		wait for 10 ns;
		t_blur_matrix_int <= (27,29,36,25,27,32,34,52,26,23,30,33,27,28,46,71,21,23,23,23,38,40,57,84,27,23,28,30,41,44,67,87,22,23,22,33,40,51,71,88,20,20,21,40,41,53,73,90,20,22,28,41,51,64,79,92,21,26,38,45,54,67,84,88);
		wait for 10 ns;
		t_blur_matrix_int <= (69,78,86,88,83,55,13,33,82,87,88,90,85,56,14,42,83,89,90,86,84,45,16,53,90,91,87,82,75,37,15,59,91,90,86,91,79,32,16,59,89,89,88,88,78,27,20,60,88,90,93,87,71,37,31,62,90,95,94,92,59,29,39,64);
		wait for 10 ns;
		t_blur_matrix_int <= (63,74,78,93,96,94,96,95,60,75,82,96,95,97,102,99,63,76,82,88,93,93,99,103,62,74,88,87,92,96,98,101,63,74,89,95,95,97,93,99,70,81,87,90,96,97,95,100,71,84,90,91,99,99,97,97,70,88,96,92,97,100,98,103);
		wait for 10 ns;
		t_blur_matrix_int <= (102,99,97,103,101,101,99,100,103,101,102,99,99,99,103,104,103,100,105,102,102,100,99,100,102,104,102,103,104,101,102,103,102,103,108,107,99,100,102,102,106,103,111,106,105,101,106,98,102,106,108,105,103,106,102,101,107,104,107,103,103,100,105,101);
		wait for 10 ns;
		t_blur_matrix_int <= (101,102,101,107,116,113,113,116,101,101,103,109,110,112,112,112,103,104,104,103,107,108,110,113,106,105,105,104,109,111,111,113,100,102,104,106,105,106,106,107,97,98,100,103,106,107,109,111,98,98,100,102,104,104,110,110,97,98,97,101,102,103,108,111);
		wait for 10 ns;
		t_blur_matrix_int <= (114,119,122,122,126,129,131,134,116,115,120,123,124,129,131,138,115,119,116,122,128,130,133,131,112,117,119,118,126,125,127,133,112,116,116,116,123,125,131,128,109,113,116,118,121,124,128,131,109,110,119,122,120,126,127,125,112,111,115,116,121,122,122,129);
		wait for 10 ns;
		t_blur_matrix_int <= (138,144,141,147,152,156,156,160,135,138,142,142,153,157,156,161,139,136,143,142,151,156,149,162,132,137,139,140,145,154,156,162,134,137,140,145,147,149,156,158,135,133,133,139,143,148,146,150,133,134,133,140,145,147,144,152,132,130,132,135,144,146,144,152);
		wait for 10 ns;
		t_blur_matrix_int <= (164,173,173,177,182,183,187,191,164,172,173,175,181,181,186,193,166,169,173,174,181,182,184,189,164,165,173,178,182,184,185,188,159,165,173,177,177,181,185,185,162,168,171,179,179,179,186,190,160,167,169,173,176,179,184,187,160,161,164,170,178,180,181,185);
		wait for 10 ns;
		t_blur_matrix_int <= (195,197,201,200,200,205,205,209,194,197,200,199,203,205,204,206,191,197,195,198,198,204,202,207,191,197,196,198,199,201,201,204,192,196,195,197,198,201,203,203,191,194,194,197,197,201,203,203,188,191,194,194,196,198,202,203,187,191,193,194,195,198,199,201);
		wait for 10 ns;
		t_blur_matrix_int <= (207,213,214,212,102,11,6,7,206,211,214,216,155,10,4,4,207,208,212,216,196,40,6,5,206,206,209,213,206,89,4,5,205,206,209,211,214,143,5,5,206,205,205,210,213,182,26,5,206,205,207,208,209,204,60,6,204,204,204,207,207,208,113,5);
		wait for 10 ns;
		t_blur_matrix_int <= (5,75,118,117,123,127,129,127,9,89,114,123,121,138,129,130,13,95,110,120,120,137,125,129,20,107,107,121,121,138,126,124,20,104,111,117,123,132,131,123,31,104,115,122,124,132,137,124,41,105,114,124,122,128,138,126,56,105,118,123,124,130,130,131);
		wait for 10 ns;
		t_blur_matrix_int <= (128,127,127,124,128,122,125,123,124,126,126,122,128,124,122,121,127,126,123,123,123,124,120,122,126,126,126,126,124,123,120,119,125,125,125,123,123,120,121,121,122,124,123,120,120,121,122,117,127,123,124,125,125,119,120,118,124,125,123,124,122,120,118,122);
		wait for 10 ns;
		t_blur_matrix_int <= (116,123,118,115,115,113,114,110,118,117,119,119,115,114,113,113,119,123,117,119,114,109,116,112,119,121,120,117,120,114,114,112,119,121,119,120,115,115,114,112,120,119,119,120,118,115,117,107,120,119,119,122,120,115,116,109,119,119,121,120,118,118,117,113);
		wait for 10 ns;
		t_blur_matrix_int <= (107,107,110,108,107,95,106,158,106,106,109,104,101,97,110,176,109,107,103,100,96,95,125,185,108,107,101,102,95,98,141,189,110,106,108,101,98,105,146,192,110,106,104,102,99,109,149,195,106,104,102,105,104,109,160,197,108,108,108,106,104,110,164,192);
		wait for 10 ns;
		t_blur_matrix_int <= (189,202,207,203,195,196,200,208,201,211,212,208,200,200,204,210,205,213,212,206,201,203,206,209,206,212,210,205,200,201,206,212,207,210,204,199,197,202,208,213,207,210,203,196,195,202,208,212,207,209,200,195,196,202,210,212,205,210,199,193,195,202,213,213);
		wait for 10 ns;
		t_blur_matrix_int <= (212,212,209,207,202,189,159,115,213,211,211,207,198,177,139,91,213,210,208,204,191,159,118,79,210,210,205,198,178,141,105,78,212,210,204,194,161,122,96,82,210,206,198,182,139,104,89,87,209,205,194,165,121,93,83,87,208,200,185,148,107,85,80,85);
		wait for 10 ns;
		t_blur_matrix_int <= (73,59,61,61,61,62,68,70,66,64,59,59,55,60,67,74,68,62,62,58,55,64,68,78,73,71,67,63,63,65,71,82,75,69,70,63,67,65,71,80,75,72,60,66,67,73,70,79,75,72,65,67,62,69,72,80,75,71,71,60,68,70,72,74);
		wait for 10 ns;
		t_blur_matrix_int <= (83,84,83,84,68,61,57,63,79,81,82,74,66,60,56,63,84,83,77,66,65,60,62,70,88,78,72,66,61,60,66,74,82,79,73,67,62,63,67,73,79,79,68,61,59,62,72,76,78,68,62,60,56,65,74,77,70,66,56,55,56,70,76,77);
		wait for 10 ns;
		t_blur_matrix_int <= (68,77,76,75,74,71,76,71,74,74,80,73,76,78,78,68,78,74,75,78,80,74,74,58,77,79,74,73,67,70,59,60,77,75,74,73,67,63,56,53,71,80,69,74,67,60,62,54,76,70,68,69,60,61,68,65,79,62,67,69,62,65,66,66);
		wait for 10 ns;
		t_blur_matrix_int <= (7,9,9,17,36,95,136,154,13,12,12,15,35,92,132,145,11,9,10,11,33,84,128,147,20,19,13,12,25,73,125,147,17,12,13,8,23,67,117,145,13,12,9,19,19,65,119,143,14,14,8,14,19,69,120,141,11,10,11,12,19,59,107,140);
		wait for 10 ns;
		t_blur_matrix_int <= (163,164,155,131,86,28,14,37,160,161,154,134,89,24,22,38,163,162,151,134,95,37,23,35,160,161,154,133,100,48,24,41,158,162,155,137,110,59,29,37,156,154,153,136,108,60,27,38,152,156,153,135,109,60,36,38,160,167,162,149,111,58,34,39);
		wait for 10 ns;
		t_blur_matrix_int <= (75,107,127,146,152,157,157,158,76,106,128,145,154,157,160,157,71,107,125,141,152,157,158,157,70,105,124,144,153,156,155,157,68,105,127,141,152,156,154,154,66,101,123,138,150,155,154,156,65,100,123,139,148,155,157,155,63,100,123,137,152,150,155,156);
		wait for 10 ns;
		t_blur_matrix_int <= (160,160,162,159,151,138,123,111,158,159,159,159,153,140,118,121,158,157,158,157,151,136,116,127,156,157,160,156,147,137,119,119,158,158,158,158,146,137,119,112,158,158,158,156,149,141,122,102,158,156,159,155,149,138,124,100,156,158,161,159,150,138,127,102);
		wait for 10 ns;
		t_blur_matrix_int <= (115,68,27,21,22,33,18,20,117,75,28,27,23,31,16,21,122,96,27,38,18,30,20,17,134,86,30,61,25,23,15,19,142,89,36,66,30,22,17,21,134,97,39,63,30,21,21,22,116,93,43,52,37,27,19,18,97,86,51,61,40,13,19,21);
		wait for 10 ns;
		t_blur_matrix_int <= (17,19,27,23,24,27,32,40,17,19,28,18,24,35,47,41,13,26,28,24,55,62,39,27,17,26,39,60,59,31,20,22,31,55,59,35,31,24,25,22,27,30,27,28,28,25,20,28,20,24,26,27,23,19,24,31,28,33,25,29,28,21,22,28);
		wait for 10 ns;
		t_blur_matrix_int <= (27,23,31,50,44,33,25,34,19,28,27,42,40,39,39,31,23,21,28,41,35,34,35,29,19,26,41,39,42,25,27,25,20,27,44,32,45,28,30,35,20,32,34,43,43,31,30,44,26,44,30,41,31,33,39,62,37,37,37,39,28,29,44,52);
		wait for 10 ns;
		t_blur_matrix_int <= (27,24,27,43,44,21,17,14,18,24,22,30,59,19,16,22,29,30,30,27,41,30,17,19,37,35,35,24,36,56,20,30,40,44,41,26,23,44,35,28,35,30,34,33,31,41,26,16,41,24,24,23,35,23,22,14,43,26,20,16,31,27,17,15);
		wait for 10 ns;
		t_blur_matrix_int <= (20,37,16,26,79,57,16,35,30,34,14,50,57,53,62,27,31,35,19,72,44,36,76,49,26,40,44,49,37,35,58,81,17,42,83,26,23,29,36,89,16,53,70,24,15,22,49,96,17,66,31,28,24,23,64,104,22,57,17,32,43,30,43,100);
		wait for 10 ns;
		t_blur_matrix_int <= (63,43,64,76,104,91,100,108,64,66,62,76,73,102,96,89,19,84,78,76,71,108,117,98,20,21,113,151,98,124,100,94,51,24,30,65,63,98,104,100,66,47,24,29,27,29,72,125,103,49,53,30,31,18,26,96,103,102,35,40,29,15,29,48);
		wait for 10 ns;
		t_blur_matrix_int <= (81,108,116,101,20,28,84,14,72,91,114,128,72,22,89,18,60,36,70,106,124,55,75,32,76,46,42,101,101,109,95,70,55,28,31,73,101,140,119,142,88,25,27,48,66,109,165,150,110,27,34,74,70,51,119,86,60,35,28,86,91,70,92,65);
		wait for 10 ns;
		t_blur_matrix_int <= (29,23,15,28,44,31,26,48,24,15,22,37,31,36,23,41,30,12,29,35,32,20,22,35,124,13,21,33,28,27,32,32,102,15,23,28,19,18,30,27,36,19,22,28,21,22,33,33,13,23,30,25,13,20,28,25,12,22,29,17,23,24,18,25);
		wait for 10 ns;
		t_blur_matrix_int <= (34,36,62,92,38,26,21,23,31,31,23,44,37,25,20,16,39,26,26,26,35,24,22,20,33,23,27,23,27,24,17,20,22,24,23,24,19,24,18,22,22,25,24,16,19,21,18,24,19,20,15,17,17,26,24,30,26,16,12,11,19,26,38,40);
		wait for 10 ns;
		t_blur_matrix_int <= (20,30,42,53,60,72,87,88,17,37,49,53,66,75,86,90,25,34,52,55,73,72,88,85,31,48,53,59,75,81,85,91,31,44,61,69,78,84,85,93,39,47,61,76,79,80,88,95,41,53,70,74,80,82,84,92,43,62,77,78,83,82,90,92);
		wait for 10 ns;
		t_blur_matrix_int <= (92,94,95,93,59,22,51,70,90,97,96,83,47,24,57,77,94,93,93,78,34,30,58,72,92,91,86,67,29,44,65,76,90,88,84,50,22,52,66,85,89,88,73,31,30,61,68,90,88,87,57,27,37,59,81,95,90,79,36,24,47,64,89,102);
		wait for 10 ns;
		t_blur_matrix_int <= (77,95,97,95,98,99,102,103,81,95,95,94,102,103,104,102,84,96,98,97,105,107,105,106,91,94,102,102,104,107,106,104,93,97,100,103,103,110,110,106,94,101,97,103,104,104,105,107,97,103,101,104,103,104,105,102,100,98,99,102,104,108,107,111);
		wait for 10 ns;
		t_blur_matrix_int <= (107,103,103,102,107,106,105,98,101,109,108,107,109,108,105,102,103,106,106,106,108,103,105,102,108,112,105,102,103,102,103,102,109,112,109,107,104,105,105,104,103,112,115,108,105,104,106,107,109,109,108,111,105,106,107,108,108,110,108,110,109,106,106,109);
		wait for 10 ns;
		t_blur_matrix_int <= (99,99,100,102,107,105,107,105,99,102,99,102,104,106,103,108,102,104,99,103,106,102,102,105,104,99,105,102,101,100,102,106,103,99,102,99,99,101,99,108,107,104,102,100,103,107,101,107,106,106,101,103,103,103,109,103,102,103,99,103,104,99,102,104);
		wait for 10 ns;
		t_blur_matrix_int <= (108,108,114,116,115,120,123,131,109,111,112,115,118,120,125,125,108,108,115,116,116,116,118,128,108,110,111,115,117,122,123,124,111,107,112,115,114,118,119,123,108,108,112,114,118,119,119,121,110,111,112,112,119,118,117,121,106,107,112,114,116,119,117,123);
		wait for 10 ns;
		t_blur_matrix_int <= (132,131,134,139,143,145,147,154,127,129,135,139,141,143,145,146,126,130,130,137,141,144,143,143,124,129,132,133,136,138,140,147,125,125,128,131,132,140,137,143,122,123,128,130,133,135,138,143,123,126,124,131,135,136,139,144,124,126,124,126,135,137,137,140);
		wait for 10 ns;
		t_blur_matrix_int <= (153,157,166,171,178,180,181,184,153,158,165,169,172,181,181,182,150,155,165,166,173,177,182,181,151,151,157,161,173,171,180,179,149,156,158,168,169,171,175,180,147,153,157,162,166,168,174,180,147,152,152,158,163,169,174,178,146,149,150,151,162,165,175,175);
		wait for 10 ns;
		t_blur_matrix_int <= (186,189,192,197,198,197,199,199,187,189,190,193,195,197,197,200,188,187,189,194,195,197,196,199,185,188,188,191,195,196,195,201,183,187,188,189,193,197,199,201,184,184,189,191,192,196,199,199,181,183,188,191,192,193,196,200,178,181,183,190,193,196,198,199);
		wait for 10 ns;
		t_blur_matrix_int <= (203,203,204,203,207,210,159,10,202,204,205,202,206,207,192,32,200,205,202,205,203,208,203,86,202,202,203,203,205,204,205,139,203,202,203,203,202,204,208,181,200,201,204,204,204,203,206,203,199,202,201,204,203,203,207,208,201,205,202,206,204,204,207,211);
		wait for 10 ns;
		t_blur_matrix_int <= (62,98,120,123,127,130,130,130,66,101,119,127,128,133,130,127,72,105,122,123,119,132,129,124,76,112,120,117,104,114,118,119,86,118,118,100,88,99,102,104,116,118,105,79,68,84,79,89,151,107,76,63,51,72,59,68,186,90,54,49,39,53,43,56);
		wait for 10 ns;
		t_blur_matrix_int <= (121,124,123,125,122,120,120,122,125,124,124,125,126,121,123,122,125,125,126,124,121,128,125,124,123,123,124,129,130,126,126,124,110,113,114,119,127,126,128,128,92,101,103,110,112,119,121,123,73,79,88,97,99,105,108,118,55,68,68,70,79,82,93,97);
		wait for 10 ns;
		t_blur_matrix_int <= (118,121,119,120,120,118,114,109,119,121,122,119,118,116,115,110,124,122,121,121,121,118,118,114,124,124,121,124,121,119,117,110,125,129,126,127,124,123,121,116,128,129,127,124,125,124,122,118,116,120,121,119,122,125,124,121,98,105,108,112,112,116,120,125);
		wait for 10 ns;
		t_blur_matrix_int <= (110,107,108,107,101,111,151,185,108,112,114,106,108,108,133,168,109,114,110,112,110,109,116,133,115,114,115,115,115,113,117,116,121,114,121,120,121,119,114,113,119,124,124,129,123,119,117,115,118,123,133,131,125,120,118,112,129,131,133,136,122,115,105,105);
		wait for 10 ns;
		t_blur_matrix_int <= (199,205,198,191,194,203,212,212,191,192,191,190,195,205,215,211,163,173,173,182,194,208,213,211,127,142,147,173,197,208,215,207,105,113,131,174,201,214,214,209,107,118,133,183,203,217,214,207,111,116,143,189,207,215,212,203,109,125,164,196,209,216,210,197);
		wait for 10 ns;
		t_blur_matrix_int <= (207,196,177,134,92,86,84,81,206,194,168,123,87,84,80,78,202,192,159,114,84,79,75,76,201,188,151,104,82,76,76,68,198,178,137,98,79,78,74,61,195,166,122,91,78,77,71,67,188,151,110,81,75,68,61,58,178,137,98,82,68,60,49,47);
		wait for 10 ns;
		t_blur_matrix_int <= (79,72,68,61,59,68,69,73,74,75,68,65,61,67,74,59,70,67,60,60,64,72,65,54,67,61,55,65,71,63,62,49,65,57,60,64,65,62,51,43,60,54,63,70,65,49,49,48,54,60,66,67,55,43,45,56,53,62,68,62,45,40,49,58);
		wait for 10 ns;
		t_blur_matrix_int <= (62,54,56,59,67,71,78,77,50,44,58,71,74,76,71,73,38,48,64,77,74,71,73,67,46,57,71,83,75,71,70,62,53,62,75,80,72,67,63,62,60,67,76,73,71,69,65,59,70,76,73,67,69,67,57,65,77,72,68,67,70,68,62,65);
		wait for 10 ns;
		t_blur_matrix_int <= (74,66,73,67,64,64,70,72,66,66,70,69,66,65,70,72,63,66,66,66,68,72,72,67,59,65,69,71,66,72,72,55,62,63,70,70,68,77,63,47,64,68,72,68,68,66,57,39,69,75,73,67,69,57,43,30,78,80,69,69,62,53,37,32);
		wait for 10 ns;
		t_blur_matrix_int <= (11,13,8,10,19,44,102,151,7,9,9,13,17,35,106,148,15,14,9,5,13,35,108,143,16,13,11,14,12,33,104,146,23,22,24,28,29,39,101,145,26,43,45,44,40,51,92,138,53,61,58,55,57,67,94,132,66,68,62,62,69,73,100,131);
		wait for 10 ns;
		t_blur_matrix_int <= (163,166,165,150,121,71,33,32,159,169,166,155,126,87,28,37,160,167,165,155,134,98,34,37,157,169,171,156,141,105,36,35,161,171,171,162,151,107,43,39,163,172,175,171,155,104,52,39,159,174,178,169,153,115,63,45,158,171,175,171,158,123,73,51);
		wait for 10 ns;
		t_blur_matrix_int <= (61,96,118,135,148,151,156,153,60,95,117,134,146,152,151,158,62,92,119,136,146,151,154,156,60,94,119,137,145,151,156,155,62,96,119,135,146,152,158,156,66,92,117,131,146,153,159,157,63,91,117,135,147,155,157,159,66,92,117,134,145,153,159,158);
		wait for 10 ns;
		t_blur_matrix_int <= (157,158,160,159,152,142,128,107,157,155,157,159,151,140,126,112,159,154,161,161,155,140,129,106,157,156,161,161,153,145,132,91,155,157,165,163,154,146,132,87,153,158,162,163,155,144,131,77,154,157,166,165,153,149,124,76,156,158,165,167,157,146,122,84);
		wait for 10 ns;
		t_blur_matrix_int <= (95,80,51,59,50,16,18,23,88,85,53,60,53,16,19,30,62,96,58,65,50,13,19,27,49,97,62,57,45,14,28,26,57,106,53,39,30,16,32,19,63,115,62,35,29,15,30,17,68,112,70,33,22,19,27,24,76,101,65,44,16,17,22,35);
		wait for 10 ns;
		t_blur_matrix_int <= (37,23,16,23,22,21,27,39,29,21,21,21,22,24,26,49,17,23,20,18,22,29,45,38,17,20,16,16,27,54,32,32,18,25,18,27,35,38,26,35,22,27,36,30,20,24,28,35,29,51,36,21,24,19,27,33,30,31,25,23,26,22,24,23);
		wait for 10 ns;
		t_blur_matrix_int <= (43,26,42,39,28,29,39,38,28,26,45,30,29,31,43,40,25,27,47,31,27,28,41,40,17,23,52,28,23,31,43,33,28,27,41,27,21,35,48,33,18,24,27,36,21,39,43,37,29,29,27,35,28,44,31,40,23,28,24,28,37,39,22,42);
		wait for 10 ns;
		t_blur_matrix_int <= (46,29,25,20,19,16,26,18,40,30,27,23,24,22,26,30,42,33,41,27,17,19,26,27,44,39,37,31,28,19,30,22,37,36,33,23,35,34,27,19,32,32,33,34,29,29,16,20,40,38,39,31,25,24,22,21,43,42,38,35,21,24,21,20);
		wait for 10 ns;
		t_blur_matrix_int <= (25,27,26,44,48,87,77,77,24,19,38,68,14,65,90,68,29,28,30,31,11,26,71,57,33,33,20,18,28,25,22,73,18,34,35,25,29,23,12,30,14,20,44,24,23,38,22,21,21,17,20,35,28,54,32,23,31,28,15,33,43,42,32,28);
		wait for 10 ns;
		t_blur_matrix_int <= (112,133,59,25,48,48,23,35,104,105,142,62,36,38,39,49,90,98,127,126,96,32,53,75,76,103,113,112,130,82,103,71,70,86,125,132,89,119,90,70,22,60,96,141,127,113,108,56,18,19,55,110,112,130,121,83,20,25,44,57,98,125,152,115);
		wait for 10 ns;
		t_blur_matrix_int <= (33,22,37,97,47,74,98,31,56,48,68,133,22,33,51,28,92,92,36,35,23,22,22,28,66,83,70,26,20,16,22,28,65,47,83,52,15,16,22,28,78,97,110,57,17,14,26,24,89,62,82,95,20,23,28,20,67,71,105,95,25,26,21,19);
		wait for 10 ns;
		t_blur_matrix_int <= (17,25,23,13,21,25,22,24,20,21,18,12,31,20,17,21,35,28,19,20,26,19,17,19,29,20,19,21,20,16,11,16,18,21,23,29,28,19,20,14,13,20,16,13,18,16,14,16,20,19,17,14,18,14,14,21,18,18,22,19,18,14,9,15);
		wait for 10 ns;
		t_blur_matrix_int <= (17,16,14,15,21,25,43,44,21,18,16,15,31,28,46,49,13,18,19,18,27,31,51,52,14,14,14,19,32,39,59,60,11,16,12,22,36,45,59,68,13,17,21,34,42,51,63,72,17,13,28,49,46,59,70,81,17,19,40,45,45,62,75,81);
		wait for 10 ns;
		t_blur_matrix_int <= (53,70,80,82,82,78,87,86,60,75,82,88,83,83,82,86,67,81,85,86,81,88,84,80,71,82,79,84,84,84,85,52,75,78,80,85,83,85,65,23,78,78,84,79,88,76,30,17,84,80,87,85,79,38,17,16,83,82,87,80,37,12,24,36);
		wait for 10 ns;
		t_blur_matrix_int <= (85,56,15,36,58,71,95,96,75,25,16,48,66,87,96,100,42,14,22,59,80,92,98,100,14,13,44,67,86,97,99,101,12,26,59,83,94,95,100,102,20,48,74,92,94,96,102,102,32,62,86,96,93,100,100,99,56,80,93,93,94,103,100,100);
		wait for 10 ns;
		t_blur_matrix_int <= (98,100,101,101,103,110,109,111,96,103,97,97,101,105,106,107,100,98,100,100,101,106,107,106,103,98,101,104,104,105,105,105,103,100,102,105,103,107,103,104,102,100,105,99,100,104,104,104,99,104,108,103,107,103,106,104,99,103,108,107,105,103,103,106);
		wait for 10 ns;
		t_blur_matrix_int <= (110,116,107,103,106,110,109,108,106,111,108,103,105,112,105,102,105,112,106,104,106,110,110,105,104,105,107,108,110,109,109,104,102,107,105,110,107,114,104,110,103,107,108,113,108,111,109,107,106,105,103,111,108,111,110,111,102,105,103,111,108,108,109,110);
		wait for 10 ns;
		t_blur_matrix_int <= (108,104,100,100,103,100,102,103,106,103,101,103,101,101,102,101,107,103,102,103,104,99,97,102,107,103,104,107,103,102,100,103,110,106,107,103,103,102,102,100,106,105,105,105,101,102,103,99,108,111,109,104,104,103,103,104,109,109,106,103,105,110,104,102);
		wait for 10 ns;
		t_blur_matrix_int <= (108,105,112,111,113,113,117,121,103,108,111,109,110,116,114,118,99,105,109,107,113,108,113,120,104,106,106,103,113,113,112,114,103,106,104,102,107,111,111,117,104,110,102,106,104,110,106,112,103,105,105,105,105,105,106,113,101,104,104,108,106,103,108,112);
		wait for 10 ns;
		t_blur_matrix_int <= (121,123,129,129,131,134,136,142,117,122,124,128,129,134,136,138,118,121,123,123,129,133,133,138,121,119,121,123,126,128,132,133,121,122,123,127,128,129,130,134,117,115,120,124,124,128,131,130,114,116,114,119,128,128,132,126,112,117,114,119,124,125,128,127);
		wait for 10 ns;
		t_blur_matrix_int <= (146,146,150,152,156,164,174,173,145,150,150,151,152,162,173,171,141,146,148,148,151,160,167,170,139,141,146,146,155,159,164,170,135,140,141,148,153,159,159,165,133,139,143,146,156,158,158,168,130,136,140,144,152,152,153,164,130,136,137,147,149,147,154,157);
		wait for 10 ns;
		t_blur_matrix_int <= (177,179,183,190,193,195,197,198,178,179,184,189,190,193,196,197,174,178,183,188,190,193,196,197,174,175,182,188,187,191,196,195,169,172,179,185,187,190,193,195,171,174,180,185,184,187,193,194,164,172,177,182,186,187,189,192,165,173,176,180,185,186,190,194);
		wait for 10 ns;
		t_blur_matrix_int <= (201,203,201,203,203,209,208,211,199,201,202,204,203,207,208,210,199,200,203,201,203,205,210,207,199,198,200,205,202,203,206,208,196,198,199,203,201,205,207,206,198,198,198,202,202,204,205,206,195,197,200,197,202,201,206,204,196,198,197,199,199,203,203,203);
		wait for 10 ns;
		t_blur_matrix_int <= (201,85,43,52,49,58,40,42,210,113,47,59,55,63,50,53,211,149,44,56,61,66,68,62,211,186,54,58,66,71,69,67,208,206,93,52,69,72,78,75,208,208,136,57,66,73,81,78,206,211,173,60,61,74,72,80,207,209,198,76,55,67,80,84);
		wait for 10 ns;
		t_blur_matrix_int <= (44,47,56,57,64,67,68,76,51,49,54,47,49,52,50,52,54,54,56,48,41,44,38,39,66,66,58,57,55,45,45,37,75,70,65,62,59,50,45,40,78,77,75,70,64,62,54,51,78,81,81,74,69,69,63,61,80,82,78,76,69,71,60,65);
		wait for 10 ns;
		t_blur_matrix_int <= (74,81,91,93,95,102,114,116,57,60,66,69,73,79,91,103,43,41,42,45,47,46,64,77,32,27,29,24,22,27,33,42,39,30,27,22,17,20,14,25,49,32,30,24,19,17,11,16,55,46,32,31,17,22,18,13,57,49,49,37,34,21,17,15);
		wait for 10 ns;
		t_blur_matrix_int <= (124,135,144,140,128,118,101,105,114,126,136,137,124,130,136,127,95,108,114,123,140,155,149,131,63,78,86,131,173,180,168,137,31,58,107,164,190,185,173,149,19,58,141,187,196,195,164,130,14,60,153,192,200,194,149,134,17,59,146,186,195,190,155,151);
		wait for 10 ns;
		t_blur_matrix_int <= (107,135,181,203,213,215,205,191,123,141,186,209,214,212,200,176,133,162,195,209,214,208,191,153,140,173,198,208,211,202,183,142,146,180,200,208,208,198,170,122,153,189,205,210,204,187,148,91,170,195,203,204,195,167,111,47,178,192,198,192,173,121,57,27);
		wait for 10 ns;
		t_blur_matrix_int <= (157,116,89,70,58,52,43,50,132,100,74,59,49,41,44,51,116,82,59,44,31,29,40,50,97,62,47,35,24,32,49,53,76,46,39,28,31,40,48,53,52,33,27,32,37,47,53,49,33,27,27,34,41,47,47,43,25,27,34,38,48,37,38,40);
		wait for 10 ns;
		t_blur_matrix_int <= (55,65,64,53,37,47,61,71,65,62,57,45,43,58,73,72,56,51,51,46,51,69,77,74,50,44,46,58,66,82,81,68,50,41,54,64,71,83,81,70,36,40,58,72,82,78,69,61,43,54,67,78,85,74,58,53,51,67,78,82,75,61,59,53);
		wait for 10 ns;
		t_blur_matrix_int <= (78,66,65,66,67,65,67,68,75,67,64,71,64,62,68,77,60,62,65,70,61,63,68,76,64,60,61,61,64,63,71,76,61,62,55,61,62,67,73,79,56,56,60,52,65,72,83,82,57,56,57,55,61,77,87,86,50,53,55,63,71,85,93,77);
		wait for 10 ns;
		t_blur_matrix_int <= (79,78,70,68,56,44,30,28,81,73,71,65,48,42,24,27,78,67,70,61,50,33,28,26,78,73,67,55,35,31,28,25,77,71,61,50,34,32,22,22,76,68,56,40,39,28,27,27,73,64,55,49,45,35,28,33,74,63,55,53,41,34,31,39);
		wait for 10 ns;
		t_blur_matrix_int <= (58,65,63,66,75,85,110,138,59,64,67,75,82,94,118,138,45,61,75,87,92,99,115,134,34,62,73,91,93,93,105,131,25,52,71,86,86,84,93,120,19,38,57,67,70,74,91,118,19,32,41,60,69,70,87,110,26,29,32,49,59,65,73,103);
		wait for 10 ns;
		t_blur_matrix_int <= (159,170,176,174,161,130,84,48,162,171,176,172,163,132,89,50,161,168,171,166,159,132,92,53,156,164,168,167,158,132,92,60,150,164,170,169,160,130,90,61,147,165,171,168,161,135,99,62,145,162,169,166,160,138,108,70,138,157,165,167,159,137,108,81);
		wait for 10 ns;
		t_blur_matrix_int <= (68,88,116,134,147,155,157,161,66,89,114,135,147,154,157,159,70,90,115,134,144,154,157,158,72,87,113,133,149,154,154,158,70,87,113,132,146,154,159,159,70,88,110,130,145,155,156,160,69,86,111,128,141,153,156,160,74,88,106,127,147,152,157,159);
		wait for 10 ns;
		t_blur_matrix_int <= (157,158,164,167,160,150,121,76,158,163,168,162,158,150,127,55,158,163,167,167,155,147,129,54,159,161,166,166,157,147,131,57,159,160,164,162,158,146,135,63,163,163,166,167,157,148,137,79,163,162,166,167,158,148,138,91,161,160,162,167,157,142,137,100);
		wait for 10 ns;
		t_blur_matrix_int <= (78,95,64,42,23,24,23,21,91,88,63,33,18,29,21,26,98,85,58,20,19,28,25,28,88,89,66,19,20,22,20,33,72,84,50,18,17,25,24,33,54,68,40,22,23,20,24,32,38,55,21,23,24,18,21,26,32,52,18,27,21,21,40,24);
		wait for 10 ns;
		t_blur_matrix_int <= (19,25,25,21,22,17,29,36,22,23,25,21,25,19,26,36,22,27,20,31,29,22,26,36,24,37,18,37,30,23,26,38,24,32,23,39,29,22,23,29,31,28,19,42,34,20,26,25,25,29,29,39,31,28,28,27,20,27,34,41,32,32,34,29);
		wait for 10 ns;
		t_blur_matrix_int <= (31,27,22,21,24,20,31,45,30,26,27,25,24,20,37,37,25,21,26,22,24,39,53,46,38,25,17,19,23,38,54,65,50,39,21,24,22,45,49,76,59,24,25,25,23,40,42,76,70,23,23,26,28,34,34,77,76,31,23,24,26,42,44,78);
		wait for 10 ns;
		t_blur_matrix_int <= (46,34,29,38,41,18,23,20,39,28,26,52,61,24,30,22,49,21,33,60,66,24,21,28,53,25,38,66,68,52,21,20,55,23,35,64,75,65,30,21,50,16,37,58,90,77,63,28,42,17,36,68,97,87,85,39,33,16,23,63,82,94,90,47);
		wait for 10 ns;
		t_blur_matrix_int <= (24,38,34,17,37,43,38,30,16,39,63,28,21,38,53,29,15,39,67,63,28,29,66,26,19,32,68,43,44,35,42,64,26,20,70,41,19,23,36,104,24,22,44,73,17,28,37,72,33,26,28,84,40,25,23,36,17,19,59,71,91,14,12,44);
		wait for 10 ns;
		t_blur_matrix_int <= (34,46,35,47,45,57,90,120,23,62,59,29,63,65,80,60,38,48,73,39,61,108,108,38,31,43,33,58,48,84,135,77,36,36,31,57,57,65,130,95,96,36,32,40,66,88,99,152,97,55,49,33,63,97,95,113,45,87,42,46,40,104,94,67);
		wait for 10 ns;
		t_blur_matrix_int <= (102,97,50,28,23,22,23,19,102,132,63,21,23,23,21,25,49,63,73,25,25,20,20,22,52,19,65,38,22,17,20,25,53,29,46,45,20,13,23,24,95,27,28,44,17,14,20,28,121,69,31,36,19,17,19,16,75,90,65,28,20,26,30,32);
		wait for 10 ns;
		t_blur_matrix_int <= (24,17,22,17,11,10,16,23,26,19,18,18,17,12,18,20,22,20,18,15,10,18,27,26,24,15,12,19,11,13,12,28,16,17,14,23,20,16,26,41,20,27,17,19,19,22,23,21,20,24,29,16,19,15,12,17,27,17,13,14,14,16,25,33);
		wait for 10 ns;
		t_blur_matrix_int <= (19,32,41,51,52,71,76,90,27,43,44,51,66,70,81,86,39,47,52,66,69,70,78,70,48,49,60,65,65,53,31,17,49,47,45,29,26,25,18,19,19,25,14,15,26,34,43,59,22,22,40,40,46,54,56,61,35,40,52,51,59,57,73,75);
		wait for 10 ns;
		t_blur_matrix_int <= (84,80,75,34,11,10,31,55,78,69,26,11,17,35,54,69,38,17,14,15,43,62,72,79,15,18,35,57,67,73,82,83,36,47,63,66,75,84,86,85,66,66,73,77,84,85,94,88,70,80,84,86,93,90,92,95,83,87,87,84,86,87,90,94);
		wait for 10 ns;
		t_blur_matrix_int <= (74,93,92,93,94,99,100,102,86,87,90,93,97,91,102,102,88,90,92,93,95,97,100,103,91,87,94,96,96,99,100,102,89,92,101,96,95,97,104,100,88,89,94,94,96,94,98,104,95,93,94,91,96,97,100,98,92,94,92,94,94,91,98,101);
		wait for 10 ns;
		t_blur_matrix_int <= (98,102,104,106,104,106,104,107,100,107,102,107,102,104,101,108,100,105,107,104,103,104,105,103,101,103,105,101,103,108,109,108,100,103,103,99,102,108,107,104,102,104,100,107,102,106,106,101,96,106,101,101,106,104,101,102,96,97,102,104,101,101,101,104);
		wait for 10 ns;
		t_blur_matrix_int <= (105,103,103,110,111,108,107,107,103,103,103,108,111,111,106,107,105,105,106,107,110,107,106,108,104,104,106,108,109,110,110,115,104,103,112,108,108,110,112,112,102,107,109,107,107,110,111,111,106,104,104,106,105,108,115,110,107,108,107,107,107,108,109,112);
		wait for 10 ns;
		t_blur_matrix_int <= (110,112,104,107,108,104,103,101,110,112,109,107,107,108,105,103,110,110,111,108,108,106,109,103,110,115,110,109,109,111,112,110,116,116,115,114,112,113,108,109,117,111,115,114,116,110,109,110,110,114,113,114,115,111,110,110,114,115,115,116,110,110,115,110);
		wait for 10 ns;
		t_blur_matrix_int <= (100,106,105,109,110,106,105,110,102,108,104,110,105,112,106,108,106,107,105,109,105,103,101,108,108,108,106,109,105,105,107,103,109,106,107,105,105,106,108,104,112,111,107,103,106,112,109,109,111,110,110,105,106,105,111,110,114,110,115,107,107,112,108,111);
		wait for 10 ns;
		t_blur_matrix_int <= (115,113,114,122,122,123,122,129,114,114,115,116,118,119,123,127,113,112,113,117,120,117,126,126,109,109,114,118,116,118,120,124,107,112,110,117,117,119,121,126,108,112,112,112,115,120,121,122,108,108,111,114,116,116,121,122,108,109,113,110,114,121,122,118);
		wait for 10 ns;
		t_blur_matrix_int <= (133,137,138,141,139,146,153,156,128,137,137,144,137,142,150,157,125,135,139,137,143,146,148,145,128,133,135,139,139,146,143,147,128,129,131,136,135,146,148,151,126,128,131,135,135,140,147,149,126,132,135,134,135,140,145,148,123,127,131,132,132,143,139,144);
		wait for 10 ns;
		t_blur_matrix_int <= (167,166,170,178,179,185,190,190,159,162,168,175,178,182,187,190,156,156,166,173,177,177,187,187,155,157,162,170,173,177,182,185,153,155,163,166,170,178,182,185,157,157,160,162,172,173,179,181,158,159,161,168,169,170,178,180,151,157,162,166,170,174,174,179);
		wait for 10 ns;
		t_blur_matrix_int <= (194,196,198,199,198,203,204,199,193,196,196,201,201,202,204,200,191,194,198,198,200,202,203,201,189,192,193,198,198,202,203,203,188,190,197,197,200,203,202,201,189,190,192,195,199,196,202,201,185,189,191,195,196,201,202,201,181,186,192,190,194,195,203,203);
		wait for 10 ns;
		t_blur_matrix_int <= (203,207,206,115,51,64,74,82,204,206,208,162,54,60,65,74,202,207,208,190,66,57,67,74,205,207,208,201,94,54,65,71,202,205,206,207,135,51,59,71,205,206,203,205,174,57,59,64,203,205,206,206,193,72,56,58,202,203,204,207,204,108,52,56);
		wait for 10 ns;
		t_blur_matrix_int <= (84,81,83,80,75,68,71,66,80,86,84,80,78,69,72,68,75,78,79,79,76,72,69,77,77,76,77,78,83,73,73,74,73,76,76,79,78,78,73,79,69,75,74,79,83,81,76,81,64,71,76,76,82,82,82,86,66,67,74,75,77,85,84,87);
		wait for 10 ns;
		t_blur_matrix_int <= (55,57,52,44,38,29,23,24,63,63,55,49,50,43,33,36,68,70,59,56,55,51,51,54,71,72,63,59,60,64,65,60,75,77,69,67,68,71,70,67,80,76,70,74,77,80,81,77,81,75,80,81,81,87,85,82,88,81,81,83,89,94,89,86);
		wait for 10 ns;
		t_blur_matrix_int <= (28,58,129,177,192,189,181,176,39,53,119,178,194,196,194,186,51,71,124,178,200,204,201,182,55,74,128,176,200,203,192,164,61,72,119,167,191,192,169,129,71,71,99,143,157,151,121,73,76,75,85,107,111,100,75,57,83,82,79,84,84,77,65,58);
		wait for 10 ns;
		t_blur_matrix_int <= (181,189,183,165,122,63,29,25,174,162,146,115,74,41,26,25,158,123,98,66,42,35,23,27,121,80,51,40,34,26,30,37,72,50,52,46,40,33,43,46,55,56,57,47,44,47,46,50,52,49,45,52,51,58,52,49,60,59,57,66,59,57,54,44);
		wait for 10 ns;
		t_blur_matrix_int <= (23,24,36,42,44,36,41,48,27,34,40,41,33,36,49,63,38,46,42,42,33,46,56,69,42,45,38,39,43,61,69,82,50,46,42,46,58,75,85,87,47,41,47,56,69,82,91,77,44,44,56,68,75,81,82,69,41,46,58,72,80,81,68,61);
		wait for 10 ns;
		t_blur_matrix_int <= (60,76,78,74,65,50,47,50,73,75,77,65,60,55,50,47,81,78,76,63,49,50,45,51,78,74,70,52,46,42,45,52,78,67,57,49,39,39,37,52,65,57,48,52,39,39,45,58,61,44,40,41,32,39,51,75,49,46,43,36,35,46,65,81);
		wait for 10 ns;
		t_blur_matrix_int <= (50,50,57,69,77,88,87,80,53,52,63,76,84,92,79,69,51,63,76,83,91,81,77,66,58,66,80,90,89,78,81,70,67,68,85,89,85,81,77,72,76,81,94,90,91,80,78,69,82,88,93,94,90,77,79,63,86,86,95,94,88,84,74,57);
		wait for 10 ns;
		t_blur_matrix_int <= (72,57,57,56,41,33,34,40,71,62,51,46,36,32,47,44,72,59,51,42,37,43,41,31,69,54,50,32,38,47,48,35,62,45,33,38,42,46,43,33,54,39,38,44,42,39,33,28,47,41,40,34,35,36,30,20,47,40,34,34,35,31,26,30);
		wait for 10 ns;
		t_blur_matrix_int <= (31,34,30,39,54,61,64,98,29,37,42,37,44,51,58,93,25,32,30,30,40,41,45,88,25,34,30,25,35,34,47,96,24,27,30,27,36,31,41,98,28,29,28,28,33,31,38,92,20,24,25,26,32,27,37,79,22,30,25,27,31,23,27,72);
		wait for 10 ns;
		t_blur_matrix_int <= (133,158,169,172,163,144,114,88,137,165,178,184,180,163,125,91,141,183,193,193,191,184,150,95,149,188,195,196,194,189,168,110,164,188,193,196,194,189,176,130,165,187,192,194,193,186,177,136,161,188,189,191,190,184,175,135,153,188,190,190,189,186,171,122);
		wait for 10 ns;
		t_blur_matrix_int <= (75,85,106,128,143,152,156,160,73,89,107,129,145,154,160,158,84,90,111,132,144,155,157,160,82,89,106,129,143,154,158,155,80,90,109,127,140,156,156,156,81,91,108,130,143,156,158,159,78,92,109,132,142,154,159,159,83,96,109,131,140,149,157,162);
		wait for 10 ns;
		t_blur_matrix_int <= (160,164,163,164,157,145,137,91,163,162,168,165,161,150,124,60,161,164,166,167,158,139,82,45,161,162,164,163,158,147,109,78,160,158,163,163,159,144,110,99,161,159,163,166,153,148,89,78,160,161,163,163,158,145,73,65,161,161,163,163,157,149,74,70);
		wait for 10 ns;
		t_blur_matrix_int <= (34,49,29,28,25,24,28,31,30,45,45,36,22,24,23,26,27,37,26,30,19,32,26,24,38,30,24,29,39,25,22,21,52,30,21,27,28,24,32,24,44,26,26,22,23,22,31,30,34,36,28,18,15,29,37,20,38,37,22,16,14,34,41,13);
		wait for 10 ns;
		t_blur_matrix_int <= (13,25,32,42,37,36,33,27,21,33,30,38,31,32,36,36,20,28,37,36,29,32,35,39,21,35,30,30,34,33,38,45,34,45,38,28,32,34,41,43,31,34,28,38,34,41,53,53,42,30,41,40,35,45,42,52,40,18,48,50,34,42,37,45);
		wait for 10 ns;
		t_blur_matrix_int <= (58,53,25,21,25,31,66,67,31,71,25,21,18,28,68,52,22,64,51,17,22,27,95,64,25,37,71,13,19,38,117,56,33,23,74,33,21,45,114,49,50,29,37,48,25,67,93,44,53,27,26,47,45,110,72,31,52,37,28,64,59,136,51,28);
		wait for 10 ns;
		t_blur_matrix_int <= (24,18,20,59,79,71,107,66,18,17,18,58,89,38,105,102,23,26,21,66,93,29,82,118,19,26,19,69,97,39,56,125,24,21,26,81,101,29,52,84,24,25,34,69,96,17,62,48,32,33,30,74,98,16,55,51,47,17,32,71,94,18,40,52);
		wait for 10 ns;
		t_blur_matrix_int <= (15,12,37,79,106,45,12,26,30,15,21,73,102,72,26,8,70,34,16,69,85,79,47,16,106,33,16,19,64,84,34,34,128,53,17,18,42,92,43,38,122,99,25,16,47,95,89,25,60,105,71,24,39,111,86,24,43,70,110,49,33,120,70,17);
		wait for 10 ns;
		t_blur_matrix_int <= (50,64,76,36,43,82,88,98,24,66,96,40,26,55,87,97,14,47,67,105,28,21,51,74,13,38,47,88,70,17,47,48,33,23,58,45,79,28,42,44,37,38,47,60,41,42,21,47,14,23,38,61,49,38,26,23,27,19,25,41,57,45,33,24);
		wait for 10 ns;
		t_blur_matrix_int <= (52,83,68,34,17,19,34,20,83,54,42,34,19,17,22,21,97,46,18,36,20,17,24,28,91,73,52,51,21,16,13,13,84,70,85,95,29,11,8,12,64,73,56,103,94,33,12,12,28,75,45,63,103,87,35,23,26,76,45,25,76,55,81,25);
		wait for 10 ns;
		t_blur_matrix_int <= (13,14,14,18,27,28,38,48,19,21,23,17,23,29,42,53,25,20,22,16,32,48,55,63,19,24,26,33,47,54,61,69,16,20,33,47,53,57,68,71,17,30,37,42,53,57,69,68,35,45,50,49,55,62,70,72,47,48,51,58,56,63,68,71);
		wait for 10 ns;
		t_blur_matrix_int <= (55,54,67,71,70,76,79,84,59,65,79,78,78,79,78,84,66,78,77,80,82,78,81,83,70,78,80,78,85,82,83,83,71,76,75,81,83,83,85,81,71,80,80,78,87,85,84,86,76,81,82,80,83,88,88,86,73,76,81,83,87,86,87,89);
		wait for 10 ns;
		t_blur_matrix_int <= (85,86,87,88,89,90,90,92,88,89,89,93,90,92,94,94,87,90,89,90,90,92,95,88,87,88,93,89,86,94,89,88,86,89,97,92,92,91,90,91,88,87,94,93,88,91,93,96,91,91,89,90,93,92,92,93,87,90,97,98,90,93,92,91);
		wait for 10 ns;
		t_blur_matrix_int <= (98,97,91,93,88,95,93,100,93,92,95,93,90,95,103,98,97,92,94,96,94,94,100,96,94,94,96,98,97,93,95,96,94,96,95,96,97,97,93,95,95,97,93,96,98,97,92,94,94,93,92,92,96,95,94,94,93,91,96,98,96,100,96,93);
		wait for 10 ns;
		t_blur_matrix_int <= (100,103,100,101,99,99,102,111,101,103,103,100,101,102,101,105,101,100,99,99,102,103,102,105,96,99,97,103,105,104,100,100,95,100,97,99,102,101,98,102,103,100,105,103,100,97,96,102,99,97,101,100,104,102,93,99,94,95,102,105,102,100,95,99);
		wait for 10 ns;
		t_blur_matrix_int <= (111,105,106,108,109,104,107,107,105,104,103,107,109,106,109,107,104,102,102,108,106,108,107,109,104,101,106,104,105,106,106,104,108,106,104,105,106,102,107,106,105,106,102,109,107,103,104,110,99,100,104,103,104,108,107,109,100,97,102,104,103,109,104,103);
		wait for 10 ns;
		t_blur_matrix_int <= (113,113,112,111,114,110,116,111,108,114,111,115,112,111,115,115,113,111,111,110,114,114,115,113,110,113,107,112,113,115,116,115,112,109,110,115,111,112,117,113,110,112,113,115,113,115,106,113,113,114,112,112,114,114,107,114,112,109,114,109,111,110,109,113);
		wait for 10 ns;
		t_blur_matrix_int <= (111,111,117,111,111,111,107,108,112,112,120,114,112,111,114,114,114,113,116,114,115,114,110,114,112,116,120,112,117,114,114,119,116,115,113,117,119,115,117,120,115,113,112,114,122,118,119,115,114,115,114,113,119,120,116,115,114,113,113,113,118,120,122,119);
		wait for 10 ns;
		t_blur_matrix_int <= (108,113,111,112,115,119,117,118,109,113,116,116,119,119,119,123,111,117,113,114,118,119,119,119,118,117,116,116,121,120,120,123,114,113,116,115,118,120,122,126,118,117,114,116,119,122,122,126,119,121,121,115,119,123,119,121,118,120,120,121,120,123,122,123);
		wait for 10 ns;
		t_blur_matrix_int <= (121,127,131,126,134,137,144,145,122,125,127,129,132,138,138,142,122,122,127,132,132,139,140,143,125,121,125,131,133,136,142,144,124,123,122,131,134,140,143,145,125,127,126,131,131,139,139,139,128,127,128,130,131,136,140,142,133,132,130,129,132,136,140,143);
		wait for 10 ns;
		t_blur_matrix_int <= (146,155,155,163,164,170,175,176,144,150,152,160,160,163,171,174,147,148,156,160,164,166,169,172,150,147,153,159,164,161,168,173,144,145,155,160,158,161,167,172,137,146,149,157,154,163,170,172,142,144,146,152,153,159,163,169,140,144,148,147,152,156,166,170);
		wait for 10 ns;
		t_blur_matrix_int <= (179,184,185,192,193,196,201,202,176,184,183,187,192,194,200,201,175,180,186,189,191,192,196,197,172,180,188,186,190,193,195,196,176,178,182,185,190,191,195,196,173,179,181,183,188,191,192,194,176,176,179,184,184,190,191,192,171,180,179,183,180,186,190,191);
		wait for 10 ns;
		t_blur_matrix_int <= (202,203,204,207,206,147,52,51,201,198,205,203,205,175,51,47,200,200,198,204,206,193,75,46,199,200,201,204,203,202,110,46,199,200,201,202,203,206,147,46,198,198,201,201,201,205,176,58,194,198,200,200,202,206,197,85,195,197,199,196,202,203,199,110);
		wait for 10 ns;
		t_blur_matrix_int <= (63,66,73,74,78,82,85,92,60,66,73,76,81,86,89,88,59,67,67,81,82,81,87,87,55,61,72,71,72,83,84,84,53,61,71,81,78,80,77,86,51,60,63,66,71,77,79,81,61,62,66,71,63,65,74,87,82,73,69,67,66,71,72,79);
		wait for 10 ns;
		t_blur_matrix_int <= (87,86,87,91,94,92,86,85,90,91,93,94,92,97,88,83,90,97,98,96,96,88,84,86,89,97,99,97,95,90,90,86,92,94,96,93,92,92,91,88,91,91,92,91,92,98,97,91,87,88,88,93,100,103,95,92,81,79,97,101,105,103,99,95);
		wait for 10 ns;
		t_blur_matrix_int <= (84,83,77,76,73,70,65,62,87,80,78,72,74,73,68,67,86,84,80,82,74,73,68,70,84,85,81,79,74,76,78,86,86,84,79,79,83,81,87,91,84,85,82,88,87,85,95,95,91,88,88,90,97,103,108,100,92,94,91,95,106,108,107,101);
		wait for 10 ns;
		t_blur_matrix_int <= (63,72,70,73,61,57,53,49,72,78,79,72,66,58,49,51,81,84,81,71,64,58,55,61,87,85,81,75,64,63,61,67,95,88,78,69,64,64,67,77,95,85,74,71,61,63,67,68,92,83,73,61,66,61,57,56,88,82,64,59,60,54,47,49);
		wait for 10 ns;
		t_blur_matrix_int <= (54,55,66,79,73,72,57,54,56,62,70,73,55,54,48,43,67,73,72,65,57,43,43,43,70,71,75,61,54,47,45,46,70,65,64,59,59,54,51,59,59,59,54,56,59,58,57,53,52,52,55,65,62,63,58,58,50,49,62,64,64,65,61,54);
		wait for 10 ns;
		t_blur_matrix_int <= (52,50,41,45,37,58,73,88,48,45,50,45,51,63,78,92,46,40,54,52,59,81,91,96,47,46,48,61,76,87,98,100,45,49,58,71,87,99,104,102,50,59,69,87,97,108,108,103,52,67,74,90,103,110,105,103,60,68,80,99,101,109,105,100);
		wait for 10 ns;
		t_blur_matrix_int <= (91,97,102,88,83,78,67,47,96,96,96,82,84,70,54,43,114,95,89,79,69,63,49,40,98,91,86,75,66,50,41,34,98,84,82,66,59,42,32,25,92,85,69,59,41,31,33,21,93,71,57,46,31,27,23,22,86,67,43,35,33,25,16,19);
		wait for 10 ns;
		t_blur_matrix_int <= (43,37,32,34,33,29,33,26,32,32,30,31,24,26,23,19,36,31,31,33,28,29,27,28,30,34,36,27,25,31,31,50,22,26,30,41,30,41,48,56,27,27,30,36,41,53,61,59,25,26,31,44,50,64,70,65,23,29,44,55,65,71,67,72);

	end process;

	
	write_process : process
	variable l: line;
	file outfile: text open write_mode is "C:\Modeltech_pe_edu_10.4a\examples\output.txt";
	begin
		wait until t_blur_clk = '0' and t_blur_clk'event;
		t_blur_comp0: for p in 0 to matrix_size-1 loop
			t_blur_comp1: for q in 0 to matrix_size-1 loop
				write(l, t_blur_res_matrix(p)(q));
				writeline(outfile, l);
			end loop t_blur_comp1;
		end loop t_blur_comp0;
	end process;

end tb_blur_behav;

configuration CFG_TB_top of tb_blur is
for tb_blur_behav
end for;
end CFG_TB_top;
